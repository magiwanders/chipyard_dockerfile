VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS
MACRO serv_top
  FOREIGN serv_top 0 0 ;
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  SIZE 288.885 BY 288.885 ;
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  30.94 276.64 276.8 278.24 ;
        RECT  30.94 249.44 276.8 251.04 ;
        RECT  30.94 222.24 276.8 223.84 ;
        RECT  30.94 195.04 276.8 196.64 ;
        RECT  30.94 167.84 276.8 169.44 ;
        RECT  30.94 140.64 276.8 142.24 ;
        RECT  30.94 113.44 276.8 115.04 ;
        RECT  30.94 86.24 276.8 87.84 ;
        RECT  30.94 59.04 276.8 60.64 ;
        RECT  30.94 31.84 276.8 33.44 ;
      LAYER met4 ;
        RECT  275.2 7.92 276.8 280.4 ;
        RECT  248.06 7.92 249.66 280.4 ;
        RECT  220.92 7.92 222.52 280.4 ;
        RECT  193.78 7.92 195.38 280.4 ;
        RECT  166.64 7.92 168.24 280.4 ;
        RECT  139.5 7.92 141.1 280.4 ;
        RECT  112.36 7.92 113.96 280.4 ;
        RECT  85.22 7.92 86.82 280.4 ;
        RECT  58.08 7.92 59.68 280.4 ;
        RECT  30.94 7.92 32.54 280.4 ;
      LAYER met1 ;
        RECT  4.6 279.92 284.28 280.4 ;
        RECT  4.6 274.48 284.28 274.96 ;
        RECT  4.6 269.04 284.28 269.52 ;
        RECT  4.6 263.6 284.28 264.08 ;
        RECT  4.6 258.16 284.28 258.64 ;
        RECT  4.6 252.72 284.28 253.2 ;
        RECT  4.6 247.28 284.28 247.76 ;
        RECT  4.6 241.84 284.28 242.32 ;
        RECT  4.6 236.4 284.28 236.88 ;
        RECT  4.6 230.96 284.28 231.44 ;
        RECT  4.6 225.52 284.28 226 ;
        RECT  4.6 220.08 284.28 220.56 ;
        RECT  4.6 214.64 284.28 215.12 ;
        RECT  4.6 209.2 284.28 209.68 ;
        RECT  4.6 203.76 284.28 204.24 ;
        RECT  4.6 198.32 284.28 198.8 ;
        RECT  4.6 192.88 284.28 193.36 ;
        RECT  4.6 187.44 284.28 187.92 ;
        RECT  4.6 182 284.28 182.48 ;
        RECT  4.6 176.56 284.28 177.04 ;
        RECT  4.6 171.12 284.28 171.6 ;
        RECT  4.6 165.68 284.28 166.16 ;
        RECT  4.6 160.24 284.28 160.72 ;
        RECT  4.6 154.8 284.28 155.28 ;
        RECT  4.6 149.36 284.28 149.84 ;
        RECT  4.6 143.92 284.28 144.4 ;
        RECT  4.6 138.48 284.28 138.96 ;
        RECT  4.6 133.04 284.28 133.52 ;
        RECT  4.6 127.6 284.28 128.08 ;
        RECT  4.6 122.16 284.28 122.64 ;
        RECT  4.6 116.72 284.28 117.2 ;
        RECT  4.6 111.28 284.28 111.76 ;
        RECT  4.6 105.84 284.28 106.32 ;
        RECT  4.6 100.4 284.28 100.88 ;
        RECT  4.6 94.96 284.28 95.44 ;
        RECT  4.6 89.52 284.28 90 ;
        RECT  4.6 84.08 284.28 84.56 ;
        RECT  4.6 78.64 284.28 79.12 ;
        RECT  4.6 73.2 284.28 73.68 ;
        RECT  4.6 67.76 284.28 68.24 ;
        RECT  4.6 62.32 284.28 62.8 ;
        RECT  4.6 56.88 284.28 57.36 ;
        RECT  4.6 51.44 284.28 51.92 ;
        RECT  4.6 46 284.28 46.48 ;
        RECT  4.6 40.56 284.28 41.04 ;
        RECT  4.6 35.12 284.28 35.6 ;
        RECT  4.6 29.68 284.28 30.16 ;
        RECT  4.6 24.24 284.28 24.72 ;
        RECT  4.6 18.8 284.28 19.28 ;
        RECT  4.6 13.36 284.28 13.84 ;
        RECT  4.6 7.92 284.28 8.4 ;
      VIA 276 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 276 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 276 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 276 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 276 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 276 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 276 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 276 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 276 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 276 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 248.86 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 221.72 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 194.58 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 167.44 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 140.3 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 113.16 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 86.02 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 58.88 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 277.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 250.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 223.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 195.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 168.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 141.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 114.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 87.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 59.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 31.74 32.64 via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  275.21 279.995 276.79 280.325 ;
      VIA 276 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 279.975 276.77 280.345 ;
      VIA 276 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 276 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 274.555 276.79 274.885 ;
      VIA 276 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 274.535 276.77 274.905 ;
      VIA 276 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 276 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 269.115 276.79 269.445 ;
      VIA 276 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 269.095 276.77 269.465 ;
      VIA 276 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 276 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 263.675 276.79 264.005 ;
      VIA 276 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 263.655 276.77 264.025 ;
      VIA 276 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 276 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 258.235 276.79 258.565 ;
      VIA 276 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 258.215 276.77 258.585 ;
      VIA 276 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 276 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 252.795 276.79 253.125 ;
      VIA 276 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 252.775 276.77 253.145 ;
      VIA 276 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 276 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 247.355 276.79 247.685 ;
      VIA 276 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 247.335 276.77 247.705 ;
      VIA 276 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 276 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 241.915 276.79 242.245 ;
      VIA 276 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 241.895 276.77 242.265 ;
      VIA 276 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 276 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 236.475 276.79 236.805 ;
      VIA 276 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 236.455 276.77 236.825 ;
      VIA 276 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 276 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 231.035 276.79 231.365 ;
      VIA 276 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 231.015 276.77 231.385 ;
      VIA 276 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 276 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 225.595 276.79 225.925 ;
      VIA 276 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 225.575 276.77 225.945 ;
      VIA 276 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 276 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 220.155 276.79 220.485 ;
      VIA 276 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 220.135 276.77 220.505 ;
      VIA 276 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 276 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 214.715 276.79 215.045 ;
      VIA 276 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 214.695 276.77 215.065 ;
      VIA 276 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 276 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 209.275 276.79 209.605 ;
      VIA 276 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 209.255 276.77 209.625 ;
      VIA 276 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 276 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 203.835 276.79 204.165 ;
      VIA 276 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 203.815 276.77 204.185 ;
      VIA 276 204 via3_4_1600_480_1_4_400_400 ;
      VIA 276 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 198.395 276.79 198.725 ;
      VIA 276 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 198.375 276.77 198.745 ;
      VIA 276 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 276 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 192.955 276.79 193.285 ;
      VIA 276 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 192.935 276.77 193.305 ;
      VIA 276 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 276 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 187.515 276.79 187.845 ;
      VIA 276 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 187.495 276.77 187.865 ;
      VIA 276 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 276 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 182.075 276.79 182.405 ;
      VIA 276 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 182.055 276.77 182.425 ;
      VIA 276 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 276 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 176.635 276.79 176.965 ;
      VIA 276 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 176.615 276.77 176.985 ;
      VIA 276 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 276 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 171.195 276.79 171.525 ;
      VIA 276 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 171.175 276.77 171.545 ;
      VIA 276 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 276 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 165.755 276.79 166.085 ;
      VIA 276 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 165.735 276.77 166.105 ;
      VIA 276 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 276 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 160.315 276.79 160.645 ;
      VIA 276 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 160.295 276.77 160.665 ;
      VIA 276 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 276 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 154.875 276.79 155.205 ;
      VIA 276 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 154.855 276.77 155.225 ;
      VIA 276 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 276 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 149.435 276.79 149.765 ;
      VIA 276 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 149.415 276.77 149.785 ;
      VIA 276 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 276 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 143.995 276.79 144.325 ;
      VIA 276 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 143.975 276.77 144.345 ;
      VIA 276 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 276 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 138.555 276.79 138.885 ;
      VIA 276 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 138.535 276.77 138.905 ;
      VIA 276 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 276 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 133.115 276.79 133.445 ;
      VIA 276 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 133.095 276.77 133.465 ;
      VIA 276 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 276 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 127.675 276.79 128.005 ;
      VIA 276 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 127.655 276.77 128.025 ;
      VIA 276 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 276 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 122.235 276.79 122.565 ;
      VIA 276 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 122.215 276.77 122.585 ;
      VIA 276 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 276 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 116.795 276.79 117.125 ;
      VIA 276 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 116.775 276.77 117.145 ;
      VIA 276 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 276 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 111.355 276.79 111.685 ;
      VIA 276 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 111.335 276.77 111.705 ;
      VIA 276 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 276 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 105.915 276.79 106.245 ;
      VIA 276 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 105.895 276.77 106.265 ;
      VIA 276 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 276 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 100.475 276.79 100.805 ;
      VIA 276 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 100.455 276.77 100.825 ;
      VIA 276 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 276 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 95.035 276.79 95.365 ;
      VIA 276 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 95.015 276.77 95.385 ;
      VIA 276 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 276 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 89.595 276.79 89.925 ;
      VIA 276 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 89.575 276.77 89.945 ;
      VIA 276 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 276 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 84.155 276.79 84.485 ;
      VIA 276 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 84.135 276.77 84.505 ;
      VIA 276 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 276 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 78.715 276.79 79.045 ;
      VIA 276 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 78.695 276.77 79.065 ;
      VIA 276 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 276 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 73.275 276.79 73.605 ;
      VIA 276 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 73.255 276.77 73.625 ;
      VIA 276 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 276 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 67.835 276.79 68.165 ;
      VIA 276 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 67.815 276.77 68.185 ;
      VIA 276 68 via3_4_1600_480_1_4_400_400 ;
      VIA 276 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 62.395 276.79 62.725 ;
      VIA 276 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 62.375 276.77 62.745 ;
      VIA 276 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 276 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 56.955 276.79 57.285 ;
      VIA 276 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 56.935 276.77 57.305 ;
      VIA 276 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 276 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 51.515 276.79 51.845 ;
      VIA 276 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 51.495 276.77 51.865 ;
      VIA 276 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 276 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 46.075 276.79 46.405 ;
      VIA 276 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 46.055 276.77 46.425 ;
      VIA 276 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 276 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 40.635 276.79 40.965 ;
      VIA 276 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 40.615 276.77 40.985 ;
      VIA 276 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 276 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 35.195 276.79 35.525 ;
      VIA 276 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 35.175 276.77 35.545 ;
      VIA 276 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 276 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 29.755 276.79 30.085 ;
      VIA 276 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 29.735 276.77 30.105 ;
      VIA 276 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 276 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 24.315 276.79 24.645 ;
      VIA 276 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 24.295 276.77 24.665 ;
      VIA 276 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 276 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 18.875 276.79 19.205 ;
      VIA 276 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 18.855 276.77 19.225 ;
      VIA 276 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 276 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 13.435 276.79 13.765 ;
      VIA 276 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 13.415 276.77 13.785 ;
      VIA 276 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 276 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  275.21 7.995 276.79 8.325 ;
      VIA 276 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  275.23 7.975 276.77 8.345 ;
      VIA 276 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 276 8.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 279.995 249.65 280.325 ;
      VIA 248.86 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 279.975 249.63 280.345 ;
      VIA 248.86 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 274.555 249.65 274.885 ;
      VIA 248.86 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 274.535 249.63 274.905 ;
      VIA 248.86 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 269.115 249.65 269.445 ;
      VIA 248.86 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 269.095 249.63 269.465 ;
      VIA 248.86 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 263.675 249.65 264.005 ;
      VIA 248.86 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 263.655 249.63 264.025 ;
      VIA 248.86 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 258.235 249.65 258.565 ;
      VIA 248.86 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 258.215 249.63 258.585 ;
      VIA 248.86 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 252.795 249.65 253.125 ;
      VIA 248.86 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 252.775 249.63 253.145 ;
      VIA 248.86 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 247.355 249.65 247.685 ;
      VIA 248.86 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 247.335 249.63 247.705 ;
      VIA 248.86 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 241.915 249.65 242.245 ;
      VIA 248.86 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 241.895 249.63 242.265 ;
      VIA 248.86 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 236.475 249.65 236.805 ;
      VIA 248.86 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 236.455 249.63 236.825 ;
      VIA 248.86 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 231.035 249.65 231.365 ;
      VIA 248.86 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 231.015 249.63 231.385 ;
      VIA 248.86 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 225.595 249.65 225.925 ;
      VIA 248.86 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 225.575 249.63 225.945 ;
      VIA 248.86 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 220.155 249.65 220.485 ;
      VIA 248.86 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 220.135 249.63 220.505 ;
      VIA 248.86 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 214.715 249.65 215.045 ;
      VIA 248.86 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 214.695 249.63 215.065 ;
      VIA 248.86 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 209.275 249.65 209.605 ;
      VIA 248.86 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 209.255 249.63 209.625 ;
      VIA 248.86 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 203.835 249.65 204.165 ;
      VIA 248.86 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 203.815 249.63 204.185 ;
      VIA 248.86 204 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 198.395 249.65 198.725 ;
      VIA 248.86 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 198.375 249.63 198.745 ;
      VIA 248.86 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 192.955 249.65 193.285 ;
      VIA 248.86 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 192.935 249.63 193.305 ;
      VIA 248.86 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 187.515 249.65 187.845 ;
      VIA 248.86 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 187.495 249.63 187.865 ;
      VIA 248.86 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 182.075 249.65 182.405 ;
      VIA 248.86 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 182.055 249.63 182.425 ;
      VIA 248.86 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 176.635 249.65 176.965 ;
      VIA 248.86 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 176.615 249.63 176.985 ;
      VIA 248.86 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 171.195 249.65 171.525 ;
      VIA 248.86 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 171.175 249.63 171.545 ;
      VIA 248.86 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 165.755 249.65 166.085 ;
      VIA 248.86 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 165.735 249.63 166.105 ;
      VIA 248.86 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 160.315 249.65 160.645 ;
      VIA 248.86 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 160.295 249.63 160.665 ;
      VIA 248.86 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 154.875 249.65 155.205 ;
      VIA 248.86 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 154.855 249.63 155.225 ;
      VIA 248.86 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 149.435 249.65 149.765 ;
      VIA 248.86 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 149.415 249.63 149.785 ;
      VIA 248.86 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 143.995 249.65 144.325 ;
      VIA 248.86 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 143.975 249.63 144.345 ;
      VIA 248.86 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 138.555 249.65 138.885 ;
      VIA 248.86 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 138.535 249.63 138.905 ;
      VIA 248.86 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 133.115 249.65 133.445 ;
      VIA 248.86 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 133.095 249.63 133.465 ;
      VIA 248.86 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 127.675 249.65 128.005 ;
      VIA 248.86 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 127.655 249.63 128.025 ;
      VIA 248.86 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 122.235 249.65 122.565 ;
      VIA 248.86 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 122.215 249.63 122.585 ;
      VIA 248.86 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 116.795 249.65 117.125 ;
      VIA 248.86 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 116.775 249.63 117.145 ;
      VIA 248.86 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 111.355 249.65 111.685 ;
      VIA 248.86 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 111.335 249.63 111.705 ;
      VIA 248.86 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 105.915 249.65 106.245 ;
      VIA 248.86 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 105.895 249.63 106.265 ;
      VIA 248.86 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 100.475 249.65 100.805 ;
      VIA 248.86 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 100.455 249.63 100.825 ;
      VIA 248.86 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 95.035 249.65 95.365 ;
      VIA 248.86 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 95.015 249.63 95.385 ;
      VIA 248.86 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 89.595 249.65 89.925 ;
      VIA 248.86 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 89.575 249.63 89.945 ;
      VIA 248.86 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 84.155 249.65 84.485 ;
      VIA 248.86 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 84.135 249.63 84.505 ;
      VIA 248.86 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 78.715 249.65 79.045 ;
      VIA 248.86 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 78.695 249.63 79.065 ;
      VIA 248.86 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 73.275 249.65 73.605 ;
      VIA 248.86 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 73.255 249.63 73.625 ;
      VIA 248.86 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 67.835 249.65 68.165 ;
      VIA 248.86 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 67.815 249.63 68.185 ;
      VIA 248.86 68 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 62.395 249.65 62.725 ;
      VIA 248.86 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 62.375 249.63 62.745 ;
      VIA 248.86 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 56.955 249.65 57.285 ;
      VIA 248.86 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 56.935 249.63 57.305 ;
      VIA 248.86 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 51.515 249.65 51.845 ;
      VIA 248.86 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 51.495 249.63 51.865 ;
      VIA 248.86 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 46.075 249.65 46.405 ;
      VIA 248.86 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 46.055 249.63 46.425 ;
      VIA 248.86 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 40.635 249.65 40.965 ;
      VIA 248.86 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 40.615 249.63 40.985 ;
      VIA 248.86 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 35.195 249.65 35.525 ;
      VIA 248.86 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 35.175 249.63 35.545 ;
      VIA 248.86 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 29.755 249.65 30.085 ;
      VIA 248.86 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 29.735 249.63 30.105 ;
      VIA 248.86 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 24.315 249.65 24.645 ;
      VIA 248.86 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 24.295 249.63 24.665 ;
      VIA 248.86 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 18.875 249.65 19.205 ;
      VIA 248.86 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 18.855 249.63 19.225 ;
      VIA 248.86 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 13.435 249.65 13.765 ;
      VIA 248.86 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 13.415 249.63 13.785 ;
      VIA 248.86 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  248.07 7.995 249.65 8.325 ;
      VIA 248.86 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  248.09 7.975 249.63 8.345 ;
      VIA 248.86 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 248.86 8.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 279.995 222.51 280.325 ;
      VIA 221.72 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 279.975 222.49 280.345 ;
      VIA 221.72 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 274.555 222.51 274.885 ;
      VIA 221.72 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 274.535 222.49 274.905 ;
      VIA 221.72 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 269.115 222.51 269.445 ;
      VIA 221.72 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 269.095 222.49 269.465 ;
      VIA 221.72 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 263.675 222.51 264.005 ;
      VIA 221.72 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 263.655 222.49 264.025 ;
      VIA 221.72 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 258.235 222.51 258.565 ;
      VIA 221.72 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 258.215 222.49 258.585 ;
      VIA 221.72 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 252.795 222.51 253.125 ;
      VIA 221.72 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 252.775 222.49 253.145 ;
      VIA 221.72 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 247.355 222.51 247.685 ;
      VIA 221.72 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 247.335 222.49 247.705 ;
      VIA 221.72 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 241.915 222.51 242.245 ;
      VIA 221.72 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 241.895 222.49 242.265 ;
      VIA 221.72 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 236.475 222.51 236.805 ;
      VIA 221.72 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 236.455 222.49 236.825 ;
      VIA 221.72 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 231.035 222.51 231.365 ;
      VIA 221.72 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 231.015 222.49 231.385 ;
      VIA 221.72 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 225.595 222.51 225.925 ;
      VIA 221.72 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 225.575 222.49 225.945 ;
      VIA 221.72 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 220.155 222.51 220.485 ;
      VIA 221.72 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 220.135 222.49 220.505 ;
      VIA 221.72 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 214.715 222.51 215.045 ;
      VIA 221.72 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 214.695 222.49 215.065 ;
      VIA 221.72 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 209.275 222.51 209.605 ;
      VIA 221.72 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 209.255 222.49 209.625 ;
      VIA 221.72 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 203.835 222.51 204.165 ;
      VIA 221.72 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 203.815 222.49 204.185 ;
      VIA 221.72 204 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 198.395 222.51 198.725 ;
      VIA 221.72 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 198.375 222.49 198.745 ;
      VIA 221.72 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 192.955 222.51 193.285 ;
      VIA 221.72 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 192.935 222.49 193.305 ;
      VIA 221.72 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 187.515 222.51 187.845 ;
      VIA 221.72 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 187.495 222.49 187.865 ;
      VIA 221.72 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 182.075 222.51 182.405 ;
      VIA 221.72 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 182.055 222.49 182.425 ;
      VIA 221.72 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 176.635 222.51 176.965 ;
      VIA 221.72 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 176.615 222.49 176.985 ;
      VIA 221.72 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 171.195 222.51 171.525 ;
      VIA 221.72 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 171.175 222.49 171.545 ;
      VIA 221.72 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 165.755 222.51 166.085 ;
      VIA 221.72 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 165.735 222.49 166.105 ;
      VIA 221.72 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 160.315 222.51 160.645 ;
      VIA 221.72 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 160.295 222.49 160.665 ;
      VIA 221.72 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 154.875 222.51 155.205 ;
      VIA 221.72 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 154.855 222.49 155.225 ;
      VIA 221.72 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 149.435 222.51 149.765 ;
      VIA 221.72 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 149.415 222.49 149.785 ;
      VIA 221.72 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 143.995 222.51 144.325 ;
      VIA 221.72 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 143.975 222.49 144.345 ;
      VIA 221.72 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 138.555 222.51 138.885 ;
      VIA 221.72 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 138.535 222.49 138.905 ;
      VIA 221.72 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 133.115 222.51 133.445 ;
      VIA 221.72 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 133.095 222.49 133.465 ;
      VIA 221.72 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 127.675 222.51 128.005 ;
      VIA 221.72 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 127.655 222.49 128.025 ;
      VIA 221.72 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 122.235 222.51 122.565 ;
      VIA 221.72 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 122.215 222.49 122.585 ;
      VIA 221.72 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 116.795 222.51 117.125 ;
      VIA 221.72 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 116.775 222.49 117.145 ;
      VIA 221.72 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 111.355 222.51 111.685 ;
      VIA 221.72 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 111.335 222.49 111.705 ;
      VIA 221.72 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 105.915 222.51 106.245 ;
      VIA 221.72 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 105.895 222.49 106.265 ;
      VIA 221.72 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 100.475 222.51 100.805 ;
      VIA 221.72 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 100.455 222.49 100.825 ;
      VIA 221.72 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 95.035 222.51 95.365 ;
      VIA 221.72 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 95.015 222.49 95.385 ;
      VIA 221.72 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 89.595 222.51 89.925 ;
      VIA 221.72 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 89.575 222.49 89.945 ;
      VIA 221.72 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 84.155 222.51 84.485 ;
      VIA 221.72 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 84.135 222.49 84.505 ;
      VIA 221.72 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 78.715 222.51 79.045 ;
      VIA 221.72 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 78.695 222.49 79.065 ;
      VIA 221.72 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 73.275 222.51 73.605 ;
      VIA 221.72 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 73.255 222.49 73.625 ;
      VIA 221.72 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 67.835 222.51 68.165 ;
      VIA 221.72 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 67.815 222.49 68.185 ;
      VIA 221.72 68 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 62.395 222.51 62.725 ;
      VIA 221.72 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 62.375 222.49 62.745 ;
      VIA 221.72 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 56.955 222.51 57.285 ;
      VIA 221.72 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 56.935 222.49 57.305 ;
      VIA 221.72 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 51.515 222.51 51.845 ;
      VIA 221.72 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 51.495 222.49 51.865 ;
      VIA 221.72 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 46.075 222.51 46.405 ;
      VIA 221.72 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 46.055 222.49 46.425 ;
      VIA 221.72 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 40.635 222.51 40.965 ;
      VIA 221.72 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 40.615 222.49 40.985 ;
      VIA 221.72 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 35.195 222.51 35.525 ;
      VIA 221.72 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 35.175 222.49 35.545 ;
      VIA 221.72 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 29.755 222.51 30.085 ;
      VIA 221.72 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 29.735 222.49 30.105 ;
      VIA 221.72 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 24.315 222.51 24.645 ;
      VIA 221.72 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 24.295 222.49 24.665 ;
      VIA 221.72 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 18.875 222.51 19.205 ;
      VIA 221.72 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 18.855 222.49 19.225 ;
      VIA 221.72 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 13.435 222.51 13.765 ;
      VIA 221.72 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 13.415 222.49 13.785 ;
      VIA 221.72 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  220.93 7.995 222.51 8.325 ;
      VIA 221.72 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  220.95 7.975 222.49 8.345 ;
      VIA 221.72 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 221.72 8.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 279.995 195.37 280.325 ;
      VIA 194.58 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 279.975 195.35 280.345 ;
      VIA 194.58 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 274.555 195.37 274.885 ;
      VIA 194.58 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 274.535 195.35 274.905 ;
      VIA 194.58 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 269.115 195.37 269.445 ;
      VIA 194.58 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 269.095 195.35 269.465 ;
      VIA 194.58 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 263.675 195.37 264.005 ;
      VIA 194.58 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 263.655 195.35 264.025 ;
      VIA 194.58 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 258.235 195.37 258.565 ;
      VIA 194.58 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 258.215 195.35 258.585 ;
      VIA 194.58 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 252.795 195.37 253.125 ;
      VIA 194.58 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 252.775 195.35 253.145 ;
      VIA 194.58 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 247.355 195.37 247.685 ;
      VIA 194.58 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 247.335 195.35 247.705 ;
      VIA 194.58 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 241.915 195.37 242.245 ;
      VIA 194.58 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 241.895 195.35 242.265 ;
      VIA 194.58 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 236.475 195.37 236.805 ;
      VIA 194.58 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 236.455 195.35 236.825 ;
      VIA 194.58 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 231.035 195.37 231.365 ;
      VIA 194.58 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 231.015 195.35 231.385 ;
      VIA 194.58 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 225.595 195.37 225.925 ;
      VIA 194.58 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 225.575 195.35 225.945 ;
      VIA 194.58 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 220.155 195.37 220.485 ;
      VIA 194.58 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 220.135 195.35 220.505 ;
      VIA 194.58 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 214.715 195.37 215.045 ;
      VIA 194.58 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 214.695 195.35 215.065 ;
      VIA 194.58 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 209.275 195.37 209.605 ;
      VIA 194.58 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 209.255 195.35 209.625 ;
      VIA 194.58 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 203.835 195.37 204.165 ;
      VIA 194.58 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 203.815 195.35 204.185 ;
      VIA 194.58 204 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 198.395 195.37 198.725 ;
      VIA 194.58 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 198.375 195.35 198.745 ;
      VIA 194.58 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 192.955 195.37 193.285 ;
      VIA 194.58 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 192.935 195.35 193.305 ;
      VIA 194.58 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 187.515 195.37 187.845 ;
      VIA 194.58 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 187.495 195.35 187.865 ;
      VIA 194.58 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 182.075 195.37 182.405 ;
      VIA 194.58 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 182.055 195.35 182.425 ;
      VIA 194.58 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 176.635 195.37 176.965 ;
      VIA 194.58 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 176.615 195.35 176.985 ;
      VIA 194.58 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 171.195 195.37 171.525 ;
      VIA 194.58 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 171.175 195.35 171.545 ;
      VIA 194.58 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 165.755 195.37 166.085 ;
      VIA 194.58 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 165.735 195.35 166.105 ;
      VIA 194.58 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 160.315 195.37 160.645 ;
      VIA 194.58 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 160.295 195.35 160.665 ;
      VIA 194.58 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 154.875 195.37 155.205 ;
      VIA 194.58 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 154.855 195.35 155.225 ;
      VIA 194.58 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 149.435 195.37 149.765 ;
      VIA 194.58 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 149.415 195.35 149.785 ;
      VIA 194.58 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 143.995 195.37 144.325 ;
      VIA 194.58 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 143.975 195.35 144.345 ;
      VIA 194.58 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 138.555 195.37 138.885 ;
      VIA 194.58 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 138.535 195.35 138.905 ;
      VIA 194.58 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 133.115 195.37 133.445 ;
      VIA 194.58 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 133.095 195.35 133.465 ;
      VIA 194.58 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 127.675 195.37 128.005 ;
      VIA 194.58 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 127.655 195.35 128.025 ;
      VIA 194.58 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 122.235 195.37 122.565 ;
      VIA 194.58 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 122.215 195.35 122.585 ;
      VIA 194.58 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 116.795 195.37 117.125 ;
      VIA 194.58 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 116.775 195.35 117.145 ;
      VIA 194.58 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 111.355 195.37 111.685 ;
      VIA 194.58 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 111.335 195.35 111.705 ;
      VIA 194.58 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 105.915 195.37 106.245 ;
      VIA 194.58 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 105.895 195.35 106.265 ;
      VIA 194.58 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 100.475 195.37 100.805 ;
      VIA 194.58 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 100.455 195.35 100.825 ;
      VIA 194.58 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 95.035 195.37 95.365 ;
      VIA 194.58 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 95.015 195.35 95.385 ;
      VIA 194.58 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 89.595 195.37 89.925 ;
      VIA 194.58 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 89.575 195.35 89.945 ;
      VIA 194.58 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 84.155 195.37 84.485 ;
      VIA 194.58 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 84.135 195.35 84.505 ;
      VIA 194.58 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 78.715 195.37 79.045 ;
      VIA 194.58 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 78.695 195.35 79.065 ;
      VIA 194.58 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 73.275 195.37 73.605 ;
      VIA 194.58 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 73.255 195.35 73.625 ;
      VIA 194.58 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 67.835 195.37 68.165 ;
      VIA 194.58 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 67.815 195.35 68.185 ;
      VIA 194.58 68 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 62.395 195.37 62.725 ;
      VIA 194.58 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 62.375 195.35 62.745 ;
      VIA 194.58 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 56.955 195.37 57.285 ;
      VIA 194.58 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 56.935 195.35 57.305 ;
      VIA 194.58 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 51.515 195.37 51.845 ;
      VIA 194.58 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 51.495 195.35 51.865 ;
      VIA 194.58 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 46.075 195.37 46.405 ;
      VIA 194.58 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 46.055 195.35 46.425 ;
      VIA 194.58 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 40.635 195.37 40.965 ;
      VIA 194.58 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 40.615 195.35 40.985 ;
      VIA 194.58 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 35.195 195.37 35.525 ;
      VIA 194.58 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 35.175 195.35 35.545 ;
      VIA 194.58 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 29.755 195.37 30.085 ;
      VIA 194.58 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 29.735 195.35 30.105 ;
      VIA 194.58 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 24.315 195.37 24.645 ;
      VIA 194.58 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 24.295 195.35 24.665 ;
      VIA 194.58 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 18.875 195.37 19.205 ;
      VIA 194.58 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 18.855 195.35 19.225 ;
      VIA 194.58 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 13.435 195.37 13.765 ;
      VIA 194.58 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 13.415 195.35 13.785 ;
      VIA 194.58 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  193.79 7.995 195.37 8.325 ;
      VIA 194.58 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  193.81 7.975 195.35 8.345 ;
      VIA 194.58 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 194.58 8.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 279.995 168.23 280.325 ;
      VIA 167.44 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 279.975 168.21 280.345 ;
      VIA 167.44 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 274.555 168.23 274.885 ;
      VIA 167.44 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 274.535 168.21 274.905 ;
      VIA 167.44 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 269.115 168.23 269.445 ;
      VIA 167.44 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 269.095 168.21 269.465 ;
      VIA 167.44 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 263.675 168.23 264.005 ;
      VIA 167.44 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 263.655 168.21 264.025 ;
      VIA 167.44 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 258.235 168.23 258.565 ;
      VIA 167.44 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 258.215 168.21 258.585 ;
      VIA 167.44 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 252.795 168.23 253.125 ;
      VIA 167.44 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 252.775 168.21 253.145 ;
      VIA 167.44 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 247.355 168.23 247.685 ;
      VIA 167.44 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 247.335 168.21 247.705 ;
      VIA 167.44 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 241.915 168.23 242.245 ;
      VIA 167.44 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 241.895 168.21 242.265 ;
      VIA 167.44 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 236.475 168.23 236.805 ;
      VIA 167.44 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 236.455 168.21 236.825 ;
      VIA 167.44 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 231.035 168.23 231.365 ;
      VIA 167.44 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 231.015 168.21 231.385 ;
      VIA 167.44 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 225.595 168.23 225.925 ;
      VIA 167.44 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 225.575 168.21 225.945 ;
      VIA 167.44 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 220.155 168.23 220.485 ;
      VIA 167.44 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 220.135 168.21 220.505 ;
      VIA 167.44 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 214.715 168.23 215.045 ;
      VIA 167.44 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 214.695 168.21 215.065 ;
      VIA 167.44 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 209.275 168.23 209.605 ;
      VIA 167.44 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 209.255 168.21 209.625 ;
      VIA 167.44 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 203.835 168.23 204.165 ;
      VIA 167.44 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 203.815 168.21 204.185 ;
      VIA 167.44 204 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 198.395 168.23 198.725 ;
      VIA 167.44 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 198.375 168.21 198.745 ;
      VIA 167.44 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 192.955 168.23 193.285 ;
      VIA 167.44 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 192.935 168.21 193.305 ;
      VIA 167.44 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 187.515 168.23 187.845 ;
      VIA 167.44 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 187.495 168.21 187.865 ;
      VIA 167.44 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 182.075 168.23 182.405 ;
      VIA 167.44 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 182.055 168.21 182.425 ;
      VIA 167.44 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 176.635 168.23 176.965 ;
      VIA 167.44 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 176.615 168.21 176.985 ;
      VIA 167.44 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 171.195 168.23 171.525 ;
      VIA 167.44 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 171.175 168.21 171.545 ;
      VIA 167.44 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 165.755 168.23 166.085 ;
      VIA 167.44 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 165.735 168.21 166.105 ;
      VIA 167.44 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 160.315 168.23 160.645 ;
      VIA 167.44 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 160.295 168.21 160.665 ;
      VIA 167.44 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 154.875 168.23 155.205 ;
      VIA 167.44 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 154.855 168.21 155.225 ;
      VIA 167.44 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 149.435 168.23 149.765 ;
      VIA 167.44 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 149.415 168.21 149.785 ;
      VIA 167.44 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 143.995 168.23 144.325 ;
      VIA 167.44 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 143.975 168.21 144.345 ;
      VIA 167.44 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 138.555 168.23 138.885 ;
      VIA 167.44 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 138.535 168.21 138.905 ;
      VIA 167.44 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 133.115 168.23 133.445 ;
      VIA 167.44 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 133.095 168.21 133.465 ;
      VIA 167.44 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 127.675 168.23 128.005 ;
      VIA 167.44 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 127.655 168.21 128.025 ;
      VIA 167.44 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 122.235 168.23 122.565 ;
      VIA 167.44 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 122.215 168.21 122.585 ;
      VIA 167.44 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 116.795 168.23 117.125 ;
      VIA 167.44 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 116.775 168.21 117.145 ;
      VIA 167.44 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 111.355 168.23 111.685 ;
      VIA 167.44 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 111.335 168.21 111.705 ;
      VIA 167.44 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 105.915 168.23 106.245 ;
      VIA 167.44 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 105.895 168.21 106.265 ;
      VIA 167.44 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 100.475 168.23 100.805 ;
      VIA 167.44 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 100.455 168.21 100.825 ;
      VIA 167.44 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 95.035 168.23 95.365 ;
      VIA 167.44 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 95.015 168.21 95.385 ;
      VIA 167.44 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 89.595 168.23 89.925 ;
      VIA 167.44 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 89.575 168.21 89.945 ;
      VIA 167.44 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 84.155 168.23 84.485 ;
      VIA 167.44 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 84.135 168.21 84.505 ;
      VIA 167.44 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 78.715 168.23 79.045 ;
      VIA 167.44 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 78.695 168.21 79.065 ;
      VIA 167.44 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 73.275 168.23 73.605 ;
      VIA 167.44 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 73.255 168.21 73.625 ;
      VIA 167.44 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 67.835 168.23 68.165 ;
      VIA 167.44 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 67.815 168.21 68.185 ;
      VIA 167.44 68 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 62.395 168.23 62.725 ;
      VIA 167.44 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 62.375 168.21 62.745 ;
      VIA 167.44 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 56.955 168.23 57.285 ;
      VIA 167.44 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 56.935 168.21 57.305 ;
      VIA 167.44 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 51.515 168.23 51.845 ;
      VIA 167.44 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 51.495 168.21 51.865 ;
      VIA 167.44 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 46.075 168.23 46.405 ;
      VIA 167.44 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 46.055 168.21 46.425 ;
      VIA 167.44 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 40.635 168.23 40.965 ;
      VIA 167.44 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 40.615 168.21 40.985 ;
      VIA 167.44 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 35.195 168.23 35.525 ;
      VIA 167.44 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 35.175 168.21 35.545 ;
      VIA 167.44 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 29.755 168.23 30.085 ;
      VIA 167.44 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 29.735 168.21 30.105 ;
      VIA 167.44 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 24.315 168.23 24.645 ;
      VIA 167.44 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 24.295 168.21 24.665 ;
      VIA 167.44 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 18.875 168.23 19.205 ;
      VIA 167.44 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 18.855 168.21 19.225 ;
      VIA 167.44 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 13.435 168.23 13.765 ;
      VIA 167.44 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 13.415 168.21 13.785 ;
      VIA 167.44 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  166.65 7.995 168.23 8.325 ;
      VIA 167.44 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  166.67 7.975 168.21 8.345 ;
      VIA 167.44 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 167.44 8.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 279.995 141.09 280.325 ;
      VIA 140.3 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 279.975 141.07 280.345 ;
      VIA 140.3 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 274.555 141.09 274.885 ;
      VIA 140.3 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 274.535 141.07 274.905 ;
      VIA 140.3 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 269.115 141.09 269.445 ;
      VIA 140.3 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 269.095 141.07 269.465 ;
      VIA 140.3 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 263.675 141.09 264.005 ;
      VIA 140.3 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 263.655 141.07 264.025 ;
      VIA 140.3 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 258.235 141.09 258.565 ;
      VIA 140.3 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 258.215 141.07 258.585 ;
      VIA 140.3 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 252.795 141.09 253.125 ;
      VIA 140.3 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 252.775 141.07 253.145 ;
      VIA 140.3 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 247.355 141.09 247.685 ;
      VIA 140.3 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 247.335 141.07 247.705 ;
      VIA 140.3 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 241.915 141.09 242.245 ;
      VIA 140.3 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 241.895 141.07 242.265 ;
      VIA 140.3 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 236.475 141.09 236.805 ;
      VIA 140.3 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 236.455 141.07 236.825 ;
      VIA 140.3 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 231.035 141.09 231.365 ;
      VIA 140.3 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 231.015 141.07 231.385 ;
      VIA 140.3 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 225.595 141.09 225.925 ;
      VIA 140.3 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 225.575 141.07 225.945 ;
      VIA 140.3 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 220.155 141.09 220.485 ;
      VIA 140.3 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 220.135 141.07 220.505 ;
      VIA 140.3 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 214.715 141.09 215.045 ;
      VIA 140.3 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 214.695 141.07 215.065 ;
      VIA 140.3 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 209.275 141.09 209.605 ;
      VIA 140.3 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 209.255 141.07 209.625 ;
      VIA 140.3 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 203.835 141.09 204.165 ;
      VIA 140.3 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 203.815 141.07 204.185 ;
      VIA 140.3 204 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 198.395 141.09 198.725 ;
      VIA 140.3 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 198.375 141.07 198.745 ;
      VIA 140.3 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 192.955 141.09 193.285 ;
      VIA 140.3 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 192.935 141.07 193.305 ;
      VIA 140.3 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 187.515 141.09 187.845 ;
      VIA 140.3 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 187.495 141.07 187.865 ;
      VIA 140.3 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 182.075 141.09 182.405 ;
      VIA 140.3 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 182.055 141.07 182.425 ;
      VIA 140.3 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 176.635 141.09 176.965 ;
      VIA 140.3 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 176.615 141.07 176.985 ;
      VIA 140.3 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 171.195 141.09 171.525 ;
      VIA 140.3 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 171.175 141.07 171.545 ;
      VIA 140.3 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 165.755 141.09 166.085 ;
      VIA 140.3 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 165.735 141.07 166.105 ;
      VIA 140.3 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 160.315 141.09 160.645 ;
      VIA 140.3 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 160.295 141.07 160.665 ;
      VIA 140.3 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 154.875 141.09 155.205 ;
      VIA 140.3 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 154.855 141.07 155.225 ;
      VIA 140.3 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 149.435 141.09 149.765 ;
      VIA 140.3 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 149.415 141.07 149.785 ;
      VIA 140.3 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 143.995 141.09 144.325 ;
      VIA 140.3 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 143.975 141.07 144.345 ;
      VIA 140.3 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 138.555 141.09 138.885 ;
      VIA 140.3 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 138.535 141.07 138.905 ;
      VIA 140.3 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 133.115 141.09 133.445 ;
      VIA 140.3 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 133.095 141.07 133.465 ;
      VIA 140.3 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 127.675 141.09 128.005 ;
      VIA 140.3 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 127.655 141.07 128.025 ;
      VIA 140.3 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 122.235 141.09 122.565 ;
      VIA 140.3 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 122.215 141.07 122.585 ;
      VIA 140.3 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 116.795 141.09 117.125 ;
      VIA 140.3 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 116.775 141.07 117.145 ;
      VIA 140.3 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 111.355 141.09 111.685 ;
      VIA 140.3 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 111.335 141.07 111.705 ;
      VIA 140.3 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 105.915 141.09 106.245 ;
      VIA 140.3 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 105.895 141.07 106.265 ;
      VIA 140.3 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 100.475 141.09 100.805 ;
      VIA 140.3 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 100.455 141.07 100.825 ;
      VIA 140.3 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 95.035 141.09 95.365 ;
      VIA 140.3 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 95.015 141.07 95.385 ;
      VIA 140.3 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 89.595 141.09 89.925 ;
      VIA 140.3 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 89.575 141.07 89.945 ;
      VIA 140.3 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 84.155 141.09 84.485 ;
      VIA 140.3 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 84.135 141.07 84.505 ;
      VIA 140.3 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 78.715 141.09 79.045 ;
      VIA 140.3 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 78.695 141.07 79.065 ;
      VIA 140.3 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 73.275 141.09 73.605 ;
      VIA 140.3 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 73.255 141.07 73.625 ;
      VIA 140.3 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 67.835 141.09 68.165 ;
      VIA 140.3 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 67.815 141.07 68.185 ;
      VIA 140.3 68 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 62.395 141.09 62.725 ;
      VIA 140.3 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 62.375 141.07 62.745 ;
      VIA 140.3 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 56.955 141.09 57.285 ;
      VIA 140.3 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 56.935 141.07 57.305 ;
      VIA 140.3 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 51.515 141.09 51.845 ;
      VIA 140.3 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 51.495 141.07 51.865 ;
      VIA 140.3 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 46.075 141.09 46.405 ;
      VIA 140.3 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 46.055 141.07 46.425 ;
      VIA 140.3 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 40.635 141.09 40.965 ;
      VIA 140.3 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 40.615 141.07 40.985 ;
      VIA 140.3 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 35.195 141.09 35.525 ;
      VIA 140.3 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 35.175 141.07 35.545 ;
      VIA 140.3 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 29.755 141.09 30.085 ;
      VIA 140.3 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 29.735 141.07 30.105 ;
      VIA 140.3 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 24.315 141.09 24.645 ;
      VIA 140.3 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 24.295 141.07 24.665 ;
      VIA 140.3 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 18.875 141.09 19.205 ;
      VIA 140.3 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 18.855 141.07 19.225 ;
      VIA 140.3 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 13.435 141.09 13.765 ;
      VIA 140.3 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 13.415 141.07 13.785 ;
      VIA 140.3 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  139.51 7.995 141.09 8.325 ;
      VIA 140.3 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  139.53 7.975 141.07 8.345 ;
      VIA 140.3 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 140.3 8.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 279.995 113.95 280.325 ;
      VIA 113.16 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 279.975 113.93 280.345 ;
      VIA 113.16 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 274.555 113.95 274.885 ;
      VIA 113.16 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 274.535 113.93 274.905 ;
      VIA 113.16 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 269.115 113.95 269.445 ;
      VIA 113.16 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 269.095 113.93 269.465 ;
      VIA 113.16 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 263.675 113.95 264.005 ;
      VIA 113.16 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 263.655 113.93 264.025 ;
      VIA 113.16 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 258.235 113.95 258.565 ;
      VIA 113.16 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 258.215 113.93 258.585 ;
      VIA 113.16 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 252.795 113.95 253.125 ;
      VIA 113.16 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 252.775 113.93 253.145 ;
      VIA 113.16 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 247.355 113.95 247.685 ;
      VIA 113.16 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 247.335 113.93 247.705 ;
      VIA 113.16 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 241.915 113.95 242.245 ;
      VIA 113.16 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 241.895 113.93 242.265 ;
      VIA 113.16 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 236.475 113.95 236.805 ;
      VIA 113.16 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 236.455 113.93 236.825 ;
      VIA 113.16 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 231.035 113.95 231.365 ;
      VIA 113.16 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 231.015 113.93 231.385 ;
      VIA 113.16 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 225.595 113.95 225.925 ;
      VIA 113.16 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 225.575 113.93 225.945 ;
      VIA 113.16 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 220.155 113.95 220.485 ;
      VIA 113.16 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 220.135 113.93 220.505 ;
      VIA 113.16 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 214.715 113.95 215.045 ;
      VIA 113.16 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 214.695 113.93 215.065 ;
      VIA 113.16 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 209.275 113.95 209.605 ;
      VIA 113.16 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 209.255 113.93 209.625 ;
      VIA 113.16 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 203.835 113.95 204.165 ;
      VIA 113.16 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 203.815 113.93 204.185 ;
      VIA 113.16 204 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 198.395 113.95 198.725 ;
      VIA 113.16 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 198.375 113.93 198.745 ;
      VIA 113.16 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 192.955 113.95 193.285 ;
      VIA 113.16 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 192.935 113.93 193.305 ;
      VIA 113.16 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 187.515 113.95 187.845 ;
      VIA 113.16 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 187.495 113.93 187.865 ;
      VIA 113.16 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 182.075 113.95 182.405 ;
      VIA 113.16 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 182.055 113.93 182.425 ;
      VIA 113.16 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 176.635 113.95 176.965 ;
      VIA 113.16 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 176.615 113.93 176.985 ;
      VIA 113.16 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 171.195 113.95 171.525 ;
      VIA 113.16 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 171.175 113.93 171.545 ;
      VIA 113.16 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 165.755 113.95 166.085 ;
      VIA 113.16 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 165.735 113.93 166.105 ;
      VIA 113.16 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 160.315 113.95 160.645 ;
      VIA 113.16 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 160.295 113.93 160.665 ;
      VIA 113.16 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 154.875 113.95 155.205 ;
      VIA 113.16 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 154.855 113.93 155.225 ;
      VIA 113.16 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 149.435 113.95 149.765 ;
      VIA 113.16 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 149.415 113.93 149.785 ;
      VIA 113.16 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 143.995 113.95 144.325 ;
      VIA 113.16 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 143.975 113.93 144.345 ;
      VIA 113.16 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 138.555 113.95 138.885 ;
      VIA 113.16 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 138.535 113.93 138.905 ;
      VIA 113.16 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 133.115 113.95 133.445 ;
      VIA 113.16 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 133.095 113.93 133.465 ;
      VIA 113.16 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 127.675 113.95 128.005 ;
      VIA 113.16 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 127.655 113.93 128.025 ;
      VIA 113.16 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 122.235 113.95 122.565 ;
      VIA 113.16 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 122.215 113.93 122.585 ;
      VIA 113.16 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 116.795 113.95 117.125 ;
      VIA 113.16 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 116.775 113.93 117.145 ;
      VIA 113.16 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 111.355 113.95 111.685 ;
      VIA 113.16 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 111.335 113.93 111.705 ;
      VIA 113.16 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 105.915 113.95 106.245 ;
      VIA 113.16 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 105.895 113.93 106.265 ;
      VIA 113.16 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 100.475 113.95 100.805 ;
      VIA 113.16 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 100.455 113.93 100.825 ;
      VIA 113.16 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 95.035 113.95 95.365 ;
      VIA 113.16 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 95.015 113.93 95.385 ;
      VIA 113.16 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 89.595 113.95 89.925 ;
      VIA 113.16 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 89.575 113.93 89.945 ;
      VIA 113.16 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 84.155 113.95 84.485 ;
      VIA 113.16 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 84.135 113.93 84.505 ;
      VIA 113.16 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 78.715 113.95 79.045 ;
      VIA 113.16 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 78.695 113.93 79.065 ;
      VIA 113.16 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 73.275 113.95 73.605 ;
      VIA 113.16 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 73.255 113.93 73.625 ;
      VIA 113.16 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 67.835 113.95 68.165 ;
      VIA 113.16 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 67.815 113.93 68.185 ;
      VIA 113.16 68 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 62.395 113.95 62.725 ;
      VIA 113.16 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 62.375 113.93 62.745 ;
      VIA 113.16 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 56.955 113.95 57.285 ;
      VIA 113.16 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 56.935 113.93 57.305 ;
      VIA 113.16 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 51.515 113.95 51.845 ;
      VIA 113.16 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 51.495 113.93 51.865 ;
      VIA 113.16 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 46.075 113.95 46.405 ;
      VIA 113.16 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 46.055 113.93 46.425 ;
      VIA 113.16 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 40.635 113.95 40.965 ;
      VIA 113.16 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 40.615 113.93 40.985 ;
      VIA 113.16 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 35.195 113.95 35.525 ;
      VIA 113.16 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 35.175 113.93 35.545 ;
      VIA 113.16 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 29.755 113.95 30.085 ;
      VIA 113.16 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 29.735 113.93 30.105 ;
      VIA 113.16 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 24.315 113.95 24.645 ;
      VIA 113.16 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 24.295 113.93 24.665 ;
      VIA 113.16 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 18.875 113.95 19.205 ;
      VIA 113.16 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 18.855 113.93 19.225 ;
      VIA 113.16 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 13.435 113.95 13.765 ;
      VIA 113.16 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 13.415 113.93 13.785 ;
      VIA 113.16 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  112.37 7.995 113.95 8.325 ;
      VIA 113.16 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  112.39 7.975 113.93 8.345 ;
      VIA 113.16 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 113.16 8.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 279.995 86.81 280.325 ;
      VIA 86.02 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 279.975 86.79 280.345 ;
      VIA 86.02 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 274.555 86.81 274.885 ;
      VIA 86.02 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 274.535 86.79 274.905 ;
      VIA 86.02 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 269.115 86.81 269.445 ;
      VIA 86.02 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 269.095 86.79 269.465 ;
      VIA 86.02 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 263.675 86.81 264.005 ;
      VIA 86.02 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 263.655 86.79 264.025 ;
      VIA 86.02 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 258.235 86.81 258.565 ;
      VIA 86.02 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 258.215 86.79 258.585 ;
      VIA 86.02 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 252.795 86.81 253.125 ;
      VIA 86.02 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 252.775 86.79 253.145 ;
      VIA 86.02 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 247.355 86.81 247.685 ;
      VIA 86.02 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 247.335 86.79 247.705 ;
      VIA 86.02 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 241.915 86.81 242.245 ;
      VIA 86.02 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 241.895 86.79 242.265 ;
      VIA 86.02 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 236.475 86.81 236.805 ;
      VIA 86.02 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 236.455 86.79 236.825 ;
      VIA 86.02 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 231.035 86.81 231.365 ;
      VIA 86.02 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 231.015 86.79 231.385 ;
      VIA 86.02 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 225.595 86.81 225.925 ;
      VIA 86.02 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 225.575 86.79 225.945 ;
      VIA 86.02 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 220.155 86.81 220.485 ;
      VIA 86.02 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 220.135 86.79 220.505 ;
      VIA 86.02 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 214.715 86.81 215.045 ;
      VIA 86.02 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 214.695 86.79 215.065 ;
      VIA 86.02 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 209.275 86.81 209.605 ;
      VIA 86.02 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 209.255 86.79 209.625 ;
      VIA 86.02 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 203.835 86.81 204.165 ;
      VIA 86.02 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 203.815 86.79 204.185 ;
      VIA 86.02 204 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 198.395 86.81 198.725 ;
      VIA 86.02 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 198.375 86.79 198.745 ;
      VIA 86.02 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 192.955 86.81 193.285 ;
      VIA 86.02 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 192.935 86.79 193.305 ;
      VIA 86.02 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 187.515 86.81 187.845 ;
      VIA 86.02 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 187.495 86.79 187.865 ;
      VIA 86.02 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 182.075 86.81 182.405 ;
      VIA 86.02 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 182.055 86.79 182.425 ;
      VIA 86.02 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 176.635 86.81 176.965 ;
      VIA 86.02 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 176.615 86.79 176.985 ;
      VIA 86.02 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 171.195 86.81 171.525 ;
      VIA 86.02 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 171.175 86.79 171.545 ;
      VIA 86.02 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 165.755 86.81 166.085 ;
      VIA 86.02 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 165.735 86.79 166.105 ;
      VIA 86.02 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 160.315 86.81 160.645 ;
      VIA 86.02 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 160.295 86.79 160.665 ;
      VIA 86.02 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 154.875 86.81 155.205 ;
      VIA 86.02 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 154.855 86.79 155.225 ;
      VIA 86.02 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 149.435 86.81 149.765 ;
      VIA 86.02 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 149.415 86.79 149.785 ;
      VIA 86.02 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 143.995 86.81 144.325 ;
      VIA 86.02 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 143.975 86.79 144.345 ;
      VIA 86.02 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 138.555 86.81 138.885 ;
      VIA 86.02 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 138.535 86.79 138.905 ;
      VIA 86.02 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 133.115 86.81 133.445 ;
      VIA 86.02 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 133.095 86.79 133.465 ;
      VIA 86.02 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 127.675 86.81 128.005 ;
      VIA 86.02 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 127.655 86.79 128.025 ;
      VIA 86.02 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 122.235 86.81 122.565 ;
      VIA 86.02 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 122.215 86.79 122.585 ;
      VIA 86.02 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 116.795 86.81 117.125 ;
      VIA 86.02 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 116.775 86.79 117.145 ;
      VIA 86.02 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 111.355 86.81 111.685 ;
      VIA 86.02 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 111.335 86.79 111.705 ;
      VIA 86.02 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 105.915 86.81 106.245 ;
      VIA 86.02 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 105.895 86.79 106.265 ;
      VIA 86.02 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 100.475 86.81 100.805 ;
      VIA 86.02 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 100.455 86.79 100.825 ;
      VIA 86.02 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 95.035 86.81 95.365 ;
      VIA 86.02 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 95.015 86.79 95.385 ;
      VIA 86.02 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 89.595 86.81 89.925 ;
      VIA 86.02 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 89.575 86.79 89.945 ;
      VIA 86.02 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 84.155 86.81 84.485 ;
      VIA 86.02 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 84.135 86.79 84.505 ;
      VIA 86.02 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 78.715 86.81 79.045 ;
      VIA 86.02 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 78.695 86.79 79.065 ;
      VIA 86.02 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 73.275 86.81 73.605 ;
      VIA 86.02 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 73.255 86.79 73.625 ;
      VIA 86.02 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 67.835 86.81 68.165 ;
      VIA 86.02 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 67.815 86.79 68.185 ;
      VIA 86.02 68 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 62.395 86.81 62.725 ;
      VIA 86.02 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 62.375 86.79 62.745 ;
      VIA 86.02 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 56.955 86.81 57.285 ;
      VIA 86.02 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 56.935 86.79 57.305 ;
      VIA 86.02 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 51.515 86.81 51.845 ;
      VIA 86.02 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 51.495 86.79 51.865 ;
      VIA 86.02 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 46.075 86.81 46.405 ;
      VIA 86.02 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 46.055 86.79 46.425 ;
      VIA 86.02 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 40.635 86.81 40.965 ;
      VIA 86.02 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 40.615 86.79 40.985 ;
      VIA 86.02 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 35.195 86.81 35.525 ;
      VIA 86.02 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 35.175 86.79 35.545 ;
      VIA 86.02 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 29.755 86.81 30.085 ;
      VIA 86.02 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 29.735 86.79 30.105 ;
      VIA 86.02 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 24.315 86.81 24.645 ;
      VIA 86.02 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 24.295 86.79 24.665 ;
      VIA 86.02 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 18.875 86.81 19.205 ;
      VIA 86.02 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 18.855 86.79 19.225 ;
      VIA 86.02 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 13.435 86.81 13.765 ;
      VIA 86.02 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 13.415 86.79 13.785 ;
      VIA 86.02 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  85.23 7.995 86.81 8.325 ;
      VIA 86.02 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  85.25 7.975 86.79 8.345 ;
      VIA 86.02 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 86.02 8.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 279.995 59.67 280.325 ;
      VIA 58.88 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 279.975 59.65 280.345 ;
      VIA 58.88 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 274.555 59.67 274.885 ;
      VIA 58.88 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 274.535 59.65 274.905 ;
      VIA 58.88 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 269.115 59.67 269.445 ;
      VIA 58.88 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 269.095 59.65 269.465 ;
      VIA 58.88 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 263.675 59.67 264.005 ;
      VIA 58.88 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 263.655 59.65 264.025 ;
      VIA 58.88 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 258.235 59.67 258.565 ;
      VIA 58.88 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 258.215 59.65 258.585 ;
      VIA 58.88 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 252.795 59.67 253.125 ;
      VIA 58.88 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 252.775 59.65 253.145 ;
      VIA 58.88 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 247.355 59.67 247.685 ;
      VIA 58.88 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 247.335 59.65 247.705 ;
      VIA 58.88 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 241.915 59.67 242.245 ;
      VIA 58.88 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 241.895 59.65 242.265 ;
      VIA 58.88 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 236.475 59.67 236.805 ;
      VIA 58.88 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 236.455 59.65 236.825 ;
      VIA 58.88 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 231.035 59.67 231.365 ;
      VIA 58.88 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 231.015 59.65 231.385 ;
      VIA 58.88 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 225.595 59.67 225.925 ;
      VIA 58.88 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 225.575 59.65 225.945 ;
      VIA 58.88 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 220.155 59.67 220.485 ;
      VIA 58.88 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 220.135 59.65 220.505 ;
      VIA 58.88 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 214.715 59.67 215.045 ;
      VIA 58.88 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 214.695 59.65 215.065 ;
      VIA 58.88 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 209.275 59.67 209.605 ;
      VIA 58.88 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 209.255 59.65 209.625 ;
      VIA 58.88 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 203.835 59.67 204.165 ;
      VIA 58.88 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 203.815 59.65 204.185 ;
      VIA 58.88 204 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 198.395 59.67 198.725 ;
      VIA 58.88 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 198.375 59.65 198.745 ;
      VIA 58.88 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 192.955 59.67 193.285 ;
      VIA 58.88 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 192.935 59.65 193.305 ;
      VIA 58.88 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 187.515 59.67 187.845 ;
      VIA 58.88 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 187.495 59.65 187.865 ;
      VIA 58.88 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 182.075 59.67 182.405 ;
      VIA 58.88 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 182.055 59.65 182.425 ;
      VIA 58.88 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 176.635 59.67 176.965 ;
      VIA 58.88 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 176.615 59.65 176.985 ;
      VIA 58.88 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 171.195 59.67 171.525 ;
      VIA 58.88 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 171.175 59.65 171.545 ;
      VIA 58.88 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 165.755 59.67 166.085 ;
      VIA 58.88 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 165.735 59.65 166.105 ;
      VIA 58.88 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 160.315 59.67 160.645 ;
      VIA 58.88 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 160.295 59.65 160.665 ;
      VIA 58.88 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 154.875 59.67 155.205 ;
      VIA 58.88 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 154.855 59.65 155.225 ;
      VIA 58.88 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 149.435 59.67 149.765 ;
      VIA 58.88 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 149.415 59.65 149.785 ;
      VIA 58.88 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 143.995 59.67 144.325 ;
      VIA 58.88 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 143.975 59.65 144.345 ;
      VIA 58.88 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 138.555 59.67 138.885 ;
      VIA 58.88 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 138.535 59.65 138.905 ;
      VIA 58.88 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 133.115 59.67 133.445 ;
      VIA 58.88 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 133.095 59.65 133.465 ;
      VIA 58.88 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 127.675 59.67 128.005 ;
      VIA 58.88 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 127.655 59.65 128.025 ;
      VIA 58.88 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 122.235 59.67 122.565 ;
      VIA 58.88 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 122.215 59.65 122.585 ;
      VIA 58.88 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 116.795 59.67 117.125 ;
      VIA 58.88 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 116.775 59.65 117.145 ;
      VIA 58.88 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 111.355 59.67 111.685 ;
      VIA 58.88 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 111.335 59.65 111.705 ;
      VIA 58.88 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 105.915 59.67 106.245 ;
      VIA 58.88 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 105.895 59.65 106.265 ;
      VIA 58.88 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 100.475 59.67 100.805 ;
      VIA 58.88 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 100.455 59.65 100.825 ;
      VIA 58.88 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 95.035 59.67 95.365 ;
      VIA 58.88 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 95.015 59.65 95.385 ;
      VIA 58.88 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 89.595 59.67 89.925 ;
      VIA 58.88 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 89.575 59.65 89.945 ;
      VIA 58.88 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 84.155 59.67 84.485 ;
      VIA 58.88 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 84.135 59.65 84.505 ;
      VIA 58.88 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 78.715 59.67 79.045 ;
      VIA 58.88 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 78.695 59.65 79.065 ;
      VIA 58.88 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 73.275 59.67 73.605 ;
      VIA 58.88 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 73.255 59.65 73.625 ;
      VIA 58.88 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 67.835 59.67 68.165 ;
      VIA 58.88 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 67.815 59.65 68.185 ;
      VIA 58.88 68 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 62.395 59.67 62.725 ;
      VIA 58.88 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 62.375 59.65 62.745 ;
      VIA 58.88 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 56.955 59.67 57.285 ;
      VIA 58.88 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 56.935 59.65 57.305 ;
      VIA 58.88 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 51.515 59.67 51.845 ;
      VIA 58.88 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 51.495 59.65 51.865 ;
      VIA 58.88 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 46.075 59.67 46.405 ;
      VIA 58.88 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 46.055 59.65 46.425 ;
      VIA 58.88 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 40.635 59.67 40.965 ;
      VIA 58.88 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 40.615 59.65 40.985 ;
      VIA 58.88 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 35.195 59.67 35.525 ;
      VIA 58.88 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 35.175 59.65 35.545 ;
      VIA 58.88 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 29.755 59.67 30.085 ;
      VIA 58.88 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 29.735 59.65 30.105 ;
      VIA 58.88 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 24.315 59.67 24.645 ;
      VIA 58.88 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 24.295 59.65 24.665 ;
      VIA 58.88 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 18.875 59.67 19.205 ;
      VIA 58.88 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 18.855 59.65 19.225 ;
      VIA 58.88 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 13.435 59.67 13.765 ;
      VIA 58.88 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 13.415 59.65 13.785 ;
      VIA 58.88 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  58.09 7.995 59.67 8.325 ;
      VIA 58.88 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  58.11 7.975 59.65 8.345 ;
      VIA 58.88 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 58.88 8.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 279.995 32.53 280.325 ;
      VIA 31.74 280.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 279.975 32.51 280.345 ;
      VIA 31.74 280.16 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 280.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 274.555 32.53 274.885 ;
      VIA 31.74 274.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 274.535 32.51 274.905 ;
      VIA 31.74 274.72 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 274.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 269.115 32.53 269.445 ;
      VIA 31.74 269.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 269.095 32.51 269.465 ;
      VIA 31.74 269.28 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 269.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 263.675 32.53 264.005 ;
      VIA 31.74 263.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 263.655 32.51 264.025 ;
      VIA 31.74 263.84 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 263.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 258.235 32.53 258.565 ;
      VIA 31.74 258.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 258.215 32.51 258.585 ;
      VIA 31.74 258.4 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 258.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 252.795 32.53 253.125 ;
      VIA 31.74 252.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 252.775 32.51 253.145 ;
      VIA 31.74 252.96 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 252.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 247.355 32.53 247.685 ;
      VIA 31.74 247.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 247.335 32.51 247.705 ;
      VIA 31.74 247.52 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 247.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 241.915 32.53 242.245 ;
      VIA 31.74 242.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 241.895 32.51 242.265 ;
      VIA 31.74 242.08 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 242.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 236.475 32.53 236.805 ;
      VIA 31.74 236.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 236.455 32.51 236.825 ;
      VIA 31.74 236.64 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 236.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 231.035 32.53 231.365 ;
      VIA 31.74 231.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 231.015 32.51 231.385 ;
      VIA 31.74 231.2 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 231.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 225.595 32.53 225.925 ;
      VIA 31.74 225.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 225.575 32.51 225.945 ;
      VIA 31.74 225.76 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 225.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 220.155 32.53 220.485 ;
      VIA 31.74 220.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 220.135 32.51 220.505 ;
      VIA 31.74 220.32 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 220.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 214.715 32.53 215.045 ;
      VIA 31.74 214.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 214.695 32.51 215.065 ;
      VIA 31.74 214.88 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 214.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 209.275 32.53 209.605 ;
      VIA 31.74 209.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 209.255 32.51 209.625 ;
      VIA 31.74 209.44 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 209.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 203.835 32.53 204.165 ;
      VIA 31.74 204 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 203.815 32.51 204.185 ;
      VIA 31.74 204 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 204 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 198.395 32.53 198.725 ;
      VIA 31.74 198.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 198.375 32.51 198.745 ;
      VIA 31.74 198.56 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 198.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 192.955 32.53 193.285 ;
      VIA 31.74 193.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 192.935 32.51 193.305 ;
      VIA 31.74 193.12 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 193.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 187.515 32.53 187.845 ;
      VIA 31.74 187.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 187.495 32.51 187.865 ;
      VIA 31.74 187.68 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 187.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 182.075 32.53 182.405 ;
      VIA 31.74 182.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 182.055 32.51 182.425 ;
      VIA 31.74 182.24 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 182.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 176.635 32.53 176.965 ;
      VIA 31.74 176.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 176.615 32.51 176.985 ;
      VIA 31.74 176.8 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 176.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 171.195 32.53 171.525 ;
      VIA 31.74 171.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 171.175 32.51 171.545 ;
      VIA 31.74 171.36 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 171.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 165.755 32.53 166.085 ;
      VIA 31.74 165.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 165.735 32.51 166.105 ;
      VIA 31.74 165.92 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 165.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 160.315 32.53 160.645 ;
      VIA 31.74 160.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 160.295 32.51 160.665 ;
      VIA 31.74 160.48 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 160.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 154.875 32.53 155.205 ;
      VIA 31.74 155.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 154.855 32.51 155.225 ;
      VIA 31.74 155.04 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 155.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 149.435 32.53 149.765 ;
      VIA 31.74 149.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 149.415 32.51 149.785 ;
      VIA 31.74 149.6 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 149.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 143.995 32.53 144.325 ;
      VIA 31.74 144.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 143.975 32.51 144.345 ;
      VIA 31.74 144.16 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 144.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 138.555 32.53 138.885 ;
      VIA 31.74 138.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 138.535 32.51 138.905 ;
      VIA 31.74 138.72 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 138.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 133.115 32.53 133.445 ;
      VIA 31.74 133.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 133.095 32.51 133.465 ;
      VIA 31.74 133.28 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 133.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 127.675 32.53 128.005 ;
      VIA 31.74 127.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 127.655 32.51 128.025 ;
      VIA 31.74 127.84 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 127.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 122.235 32.53 122.565 ;
      VIA 31.74 122.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 122.215 32.51 122.585 ;
      VIA 31.74 122.4 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 122.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 116.795 32.53 117.125 ;
      VIA 31.74 116.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 116.775 32.51 117.145 ;
      VIA 31.74 116.96 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 116.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 111.355 32.53 111.685 ;
      VIA 31.74 111.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 111.335 32.51 111.705 ;
      VIA 31.74 111.52 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 111.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 105.915 32.53 106.245 ;
      VIA 31.74 106.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 105.895 32.51 106.265 ;
      VIA 31.74 106.08 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 106.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 100.475 32.53 100.805 ;
      VIA 31.74 100.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 100.455 32.51 100.825 ;
      VIA 31.74 100.64 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 100.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 95.035 32.53 95.365 ;
      VIA 31.74 95.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 95.015 32.51 95.385 ;
      VIA 31.74 95.2 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 95.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 89.595 32.53 89.925 ;
      VIA 31.74 89.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 89.575 32.51 89.945 ;
      VIA 31.74 89.76 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 89.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 84.155 32.53 84.485 ;
      VIA 31.74 84.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 84.135 32.51 84.505 ;
      VIA 31.74 84.32 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 84.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 78.715 32.53 79.045 ;
      VIA 31.74 78.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 78.695 32.51 79.065 ;
      VIA 31.74 78.88 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 78.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 73.275 32.53 73.605 ;
      VIA 31.74 73.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 73.255 32.51 73.625 ;
      VIA 31.74 73.44 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 73.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 67.835 32.53 68.165 ;
      VIA 31.74 68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 67.815 32.51 68.185 ;
      VIA 31.74 68 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 62.395 32.53 62.725 ;
      VIA 31.74 62.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 62.375 32.51 62.745 ;
      VIA 31.74 62.56 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 62.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 56.955 32.53 57.285 ;
      VIA 31.74 57.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 56.935 32.51 57.305 ;
      VIA 31.74 57.12 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 57.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 51.515 32.53 51.845 ;
      VIA 31.74 51.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 51.495 32.51 51.865 ;
      VIA 31.74 51.68 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 51.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 46.075 32.53 46.405 ;
      VIA 31.74 46.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 46.055 32.51 46.425 ;
      VIA 31.74 46.24 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 46.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 40.635 32.53 40.965 ;
      VIA 31.74 40.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 40.615 32.51 40.985 ;
      VIA 31.74 40.8 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 40.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 35.195 32.53 35.525 ;
      VIA 31.74 35.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 35.175 32.51 35.545 ;
      VIA 31.74 35.36 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 35.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 29.755 32.53 30.085 ;
      VIA 31.74 29.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 29.735 32.51 30.105 ;
      VIA 31.74 29.92 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 29.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 24.315 32.53 24.645 ;
      VIA 31.74 24.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 24.295 32.51 24.665 ;
      VIA 31.74 24.48 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 24.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 18.875 32.53 19.205 ;
      VIA 31.74 19.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 18.855 32.51 19.225 ;
      VIA 31.74 19.04 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 19.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 13.435 32.53 13.765 ;
      VIA 31.74 13.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 13.415 32.51 13.785 ;
      VIA 31.74 13.6 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 13.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  30.95 7.995 32.53 8.325 ;
      VIA 31.74 8.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  30.97 7.975 32.51 8.345 ;
      VIA 31.74 8.16 via3_4_1600_480_1_4_400_400 ;
      VIA 31.74 8.16 via2_3_1600_480_1_5_320_320 ;
    END
  END VDD
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER met5 ;
        RECT  17.37 263.04 263.23 264.64 ;
        RECT  17.37 235.84 263.23 237.44 ;
        RECT  17.37 208.64 263.23 210.24 ;
        RECT  17.37 181.44 263.23 183.04 ;
        RECT  17.37 154.24 263.23 155.84 ;
        RECT  17.37 127.04 263.23 128.64 ;
        RECT  17.37 99.84 263.23 101.44 ;
        RECT  17.37 72.64 263.23 74.24 ;
        RECT  17.37 45.44 263.23 47.04 ;
        RECT  17.37 18.24 263.23 19.84 ;
      LAYER met4 ;
        RECT  261.63 5.2 263.23 283.12 ;
        RECT  234.49 5.2 236.09 283.12 ;
        RECT  207.35 5.2 208.95 283.12 ;
        RECT  180.21 5.2 181.81 283.12 ;
        RECT  153.07 5.2 154.67 283.12 ;
        RECT  125.93 5.2 127.53 283.12 ;
        RECT  98.79 5.2 100.39 283.12 ;
        RECT  71.65 5.2 73.25 283.12 ;
        RECT  44.51 5.2 46.11 283.12 ;
        RECT  17.37 5.2 18.97 283.12 ;
      LAYER met1 ;
        RECT  4.6 282.64 284.28 283.12 ;
        RECT  4.6 277.2 284.28 277.68 ;
        RECT  4.6 271.76 284.28 272.24 ;
        RECT  4.6 266.32 284.28 266.8 ;
        RECT  4.6 260.88 284.28 261.36 ;
        RECT  4.6 255.44 284.28 255.92 ;
        RECT  4.6 250 284.28 250.48 ;
        RECT  4.6 244.56 284.28 245.04 ;
        RECT  4.6 239.12 284.28 239.6 ;
        RECT  4.6 233.68 284.28 234.16 ;
        RECT  4.6 228.24 284.28 228.72 ;
        RECT  4.6 222.8 284.28 223.28 ;
        RECT  4.6 217.36 284.28 217.84 ;
        RECT  4.6 211.92 284.28 212.4 ;
        RECT  4.6 206.48 284.28 206.96 ;
        RECT  4.6 201.04 284.28 201.52 ;
        RECT  4.6 195.6 284.28 196.08 ;
        RECT  4.6 190.16 284.28 190.64 ;
        RECT  4.6 184.72 284.28 185.2 ;
        RECT  4.6 179.28 284.28 179.76 ;
        RECT  4.6 173.84 284.28 174.32 ;
        RECT  4.6 168.4 284.28 168.88 ;
        RECT  4.6 162.96 284.28 163.44 ;
        RECT  4.6 157.52 284.28 158 ;
        RECT  4.6 152.08 284.28 152.56 ;
        RECT  4.6 146.64 284.28 147.12 ;
        RECT  4.6 141.2 284.28 141.68 ;
        RECT  4.6 135.76 284.28 136.24 ;
        RECT  4.6 130.32 284.28 130.8 ;
        RECT  4.6 124.88 284.28 125.36 ;
        RECT  4.6 119.44 284.28 119.92 ;
        RECT  4.6 114 284.28 114.48 ;
        RECT  4.6 108.56 284.28 109.04 ;
        RECT  4.6 103.12 284.28 103.6 ;
        RECT  4.6 97.68 284.28 98.16 ;
        RECT  4.6 92.24 284.28 92.72 ;
        RECT  4.6 86.8 284.28 87.28 ;
        RECT  4.6 81.36 284.28 81.84 ;
        RECT  4.6 75.92 284.28 76.4 ;
        RECT  4.6 70.48 284.28 70.96 ;
        RECT  4.6 65.04 284.28 65.52 ;
        RECT  4.6 59.6 284.28 60.08 ;
        RECT  4.6 54.16 284.28 54.64 ;
        RECT  4.6 48.72 284.28 49.2 ;
        RECT  4.6 43.28 284.28 43.76 ;
        RECT  4.6 37.84 284.28 38.32 ;
        RECT  4.6 32.4 284.28 32.88 ;
        RECT  4.6 26.96 284.28 27.44 ;
        RECT  4.6 21.52 284.28 22 ;
        RECT  4.6 16.08 284.28 16.56 ;
        RECT  4.6 10.64 284.28 11.12 ;
        RECT  4.6 5.2 284.28 5.68 ;
      VIA 262.43 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 262.43 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 262.43 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 262.43 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 262.43 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 262.43 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 262.43 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 262.43 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 262.43 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 262.43 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 235.29 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 208.15 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 181.01 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 153.87 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 126.73 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 99.59 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 72.45 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 45.31 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 263.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 236.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 209.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 182.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 155.04 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 127.84 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 100.64 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 73.44 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 46.24 via5_6_1600_1600_1_1_1600_1600 ;
      VIA 18.17 19.04 via5_6_1600_1600_1_1_1600_1600 ;
      LAYER met3 ;
        RECT  261.64 282.715 263.22 283.045 ;
      VIA 262.43 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 282.695 263.2 283.065 ;
      VIA 262.43 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 277.275 263.22 277.605 ;
      VIA 262.43 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 277.255 263.2 277.625 ;
      VIA 262.43 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 271.835 263.22 272.165 ;
      VIA 262.43 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 271.815 263.2 272.185 ;
      VIA 262.43 272 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 266.395 263.22 266.725 ;
      VIA 262.43 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 266.375 263.2 266.745 ;
      VIA 262.43 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 260.955 263.22 261.285 ;
      VIA 262.43 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 260.935 263.2 261.305 ;
      VIA 262.43 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 255.515 263.22 255.845 ;
      VIA 262.43 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 255.495 263.2 255.865 ;
      VIA 262.43 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 250.075 263.22 250.405 ;
      VIA 262.43 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 250.055 263.2 250.425 ;
      VIA 262.43 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 244.635 263.22 244.965 ;
      VIA 262.43 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 244.615 263.2 244.985 ;
      VIA 262.43 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 239.195 263.22 239.525 ;
      VIA 262.43 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 239.175 263.2 239.545 ;
      VIA 262.43 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 233.755 263.22 234.085 ;
      VIA 262.43 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 233.735 263.2 234.105 ;
      VIA 262.43 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 228.315 263.22 228.645 ;
      VIA 262.43 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 228.295 263.2 228.665 ;
      VIA 262.43 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 222.875 263.22 223.205 ;
      VIA 262.43 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 222.855 263.2 223.225 ;
      VIA 262.43 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 217.435 263.22 217.765 ;
      VIA 262.43 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 217.415 263.2 217.785 ;
      VIA 262.43 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 211.995 263.22 212.325 ;
      VIA 262.43 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 211.975 263.2 212.345 ;
      VIA 262.43 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 206.555 263.22 206.885 ;
      VIA 262.43 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 206.535 263.2 206.905 ;
      VIA 262.43 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 201.115 263.22 201.445 ;
      VIA 262.43 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 201.095 263.2 201.465 ;
      VIA 262.43 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 195.675 263.22 196.005 ;
      VIA 262.43 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 195.655 263.2 196.025 ;
      VIA 262.43 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 190.235 263.22 190.565 ;
      VIA 262.43 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 190.215 263.2 190.585 ;
      VIA 262.43 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 184.795 263.22 185.125 ;
      VIA 262.43 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 184.775 263.2 185.145 ;
      VIA 262.43 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 179.355 263.22 179.685 ;
      VIA 262.43 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 179.335 263.2 179.705 ;
      VIA 262.43 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 173.915 263.22 174.245 ;
      VIA 262.43 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 173.895 263.2 174.265 ;
      VIA 262.43 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 168.475 263.22 168.805 ;
      VIA 262.43 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 168.455 263.2 168.825 ;
      VIA 262.43 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 163.035 263.22 163.365 ;
      VIA 262.43 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 163.015 263.2 163.385 ;
      VIA 262.43 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 157.595 263.22 157.925 ;
      VIA 262.43 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 157.575 263.2 157.945 ;
      VIA 262.43 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 152.155 263.22 152.485 ;
      VIA 262.43 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 152.135 263.2 152.505 ;
      VIA 262.43 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 146.715 263.22 147.045 ;
      VIA 262.43 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 146.695 263.2 147.065 ;
      VIA 262.43 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 141.275 263.22 141.605 ;
      VIA 262.43 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 141.255 263.2 141.625 ;
      VIA 262.43 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 135.835 263.22 136.165 ;
      VIA 262.43 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 135.815 263.2 136.185 ;
      VIA 262.43 136 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 130.395 263.22 130.725 ;
      VIA 262.43 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 130.375 263.2 130.745 ;
      VIA 262.43 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 124.955 263.22 125.285 ;
      VIA 262.43 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 124.935 263.2 125.305 ;
      VIA 262.43 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 119.515 263.22 119.845 ;
      VIA 262.43 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 119.495 263.2 119.865 ;
      VIA 262.43 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 114.075 263.22 114.405 ;
      VIA 262.43 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 114.055 263.2 114.425 ;
      VIA 262.43 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 108.635 263.22 108.965 ;
      VIA 262.43 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 108.615 263.2 108.985 ;
      VIA 262.43 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 103.195 263.22 103.525 ;
      VIA 262.43 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 103.175 263.2 103.545 ;
      VIA 262.43 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 97.755 263.22 98.085 ;
      VIA 262.43 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 97.735 263.2 98.105 ;
      VIA 262.43 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 92.315 263.22 92.645 ;
      VIA 262.43 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 92.295 263.2 92.665 ;
      VIA 262.43 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 86.875 263.22 87.205 ;
      VIA 262.43 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 86.855 263.2 87.225 ;
      VIA 262.43 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 81.435 263.22 81.765 ;
      VIA 262.43 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 81.415 263.2 81.785 ;
      VIA 262.43 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 75.995 263.22 76.325 ;
      VIA 262.43 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 75.975 263.2 76.345 ;
      VIA 262.43 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 70.555 263.22 70.885 ;
      VIA 262.43 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 70.535 263.2 70.905 ;
      VIA 262.43 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 65.115 263.22 65.445 ;
      VIA 262.43 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 65.095 263.2 65.465 ;
      VIA 262.43 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 59.675 263.22 60.005 ;
      VIA 262.43 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 59.655 263.2 60.025 ;
      VIA 262.43 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 54.235 263.22 54.565 ;
      VIA 262.43 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 54.215 263.2 54.585 ;
      VIA 262.43 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 48.795 263.22 49.125 ;
      VIA 262.43 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 48.775 263.2 49.145 ;
      VIA 262.43 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 43.355 263.22 43.685 ;
      VIA 262.43 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 43.335 263.2 43.705 ;
      VIA 262.43 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 37.915 263.22 38.245 ;
      VIA 262.43 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 37.895 263.2 38.265 ;
      VIA 262.43 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 32.475 263.22 32.805 ;
      VIA 262.43 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 32.455 263.2 32.825 ;
      VIA 262.43 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 27.035 263.22 27.365 ;
      VIA 262.43 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 27.015 263.2 27.385 ;
      VIA 262.43 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 21.595 263.22 21.925 ;
      VIA 262.43 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 21.575 263.2 21.945 ;
      VIA 262.43 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 16.155 263.22 16.485 ;
      VIA 262.43 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 16.135 263.2 16.505 ;
      VIA 262.43 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 10.715 263.22 11.045 ;
      VIA 262.43 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 10.695 263.2 11.065 ;
      VIA 262.43 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  261.64 5.275 263.22 5.605 ;
      VIA 262.43 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  261.66 5.255 263.2 5.625 ;
      VIA 262.43 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 262.43 5.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 282.715 236.08 283.045 ;
      VIA 235.29 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 282.695 236.06 283.065 ;
      VIA 235.29 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 277.275 236.08 277.605 ;
      VIA 235.29 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 277.255 236.06 277.625 ;
      VIA 235.29 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 271.835 236.08 272.165 ;
      VIA 235.29 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 271.815 236.06 272.185 ;
      VIA 235.29 272 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 266.395 236.08 266.725 ;
      VIA 235.29 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 266.375 236.06 266.745 ;
      VIA 235.29 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 260.955 236.08 261.285 ;
      VIA 235.29 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 260.935 236.06 261.305 ;
      VIA 235.29 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 255.515 236.08 255.845 ;
      VIA 235.29 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 255.495 236.06 255.865 ;
      VIA 235.29 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 250.075 236.08 250.405 ;
      VIA 235.29 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 250.055 236.06 250.425 ;
      VIA 235.29 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 244.635 236.08 244.965 ;
      VIA 235.29 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 244.615 236.06 244.985 ;
      VIA 235.29 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 239.195 236.08 239.525 ;
      VIA 235.29 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 239.175 236.06 239.545 ;
      VIA 235.29 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 233.755 236.08 234.085 ;
      VIA 235.29 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 233.735 236.06 234.105 ;
      VIA 235.29 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 228.315 236.08 228.645 ;
      VIA 235.29 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 228.295 236.06 228.665 ;
      VIA 235.29 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 222.875 236.08 223.205 ;
      VIA 235.29 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 222.855 236.06 223.225 ;
      VIA 235.29 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 217.435 236.08 217.765 ;
      VIA 235.29 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 217.415 236.06 217.785 ;
      VIA 235.29 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 211.995 236.08 212.325 ;
      VIA 235.29 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 211.975 236.06 212.345 ;
      VIA 235.29 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 206.555 236.08 206.885 ;
      VIA 235.29 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 206.535 236.06 206.905 ;
      VIA 235.29 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 201.115 236.08 201.445 ;
      VIA 235.29 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 201.095 236.06 201.465 ;
      VIA 235.29 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 195.675 236.08 196.005 ;
      VIA 235.29 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 195.655 236.06 196.025 ;
      VIA 235.29 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 190.235 236.08 190.565 ;
      VIA 235.29 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 190.215 236.06 190.585 ;
      VIA 235.29 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 184.795 236.08 185.125 ;
      VIA 235.29 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 184.775 236.06 185.145 ;
      VIA 235.29 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 179.355 236.08 179.685 ;
      VIA 235.29 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 179.335 236.06 179.705 ;
      VIA 235.29 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 173.915 236.08 174.245 ;
      VIA 235.29 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 173.895 236.06 174.265 ;
      VIA 235.29 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 168.475 236.08 168.805 ;
      VIA 235.29 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 168.455 236.06 168.825 ;
      VIA 235.29 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 163.035 236.08 163.365 ;
      VIA 235.29 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 163.015 236.06 163.385 ;
      VIA 235.29 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 157.595 236.08 157.925 ;
      VIA 235.29 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 157.575 236.06 157.945 ;
      VIA 235.29 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 152.155 236.08 152.485 ;
      VIA 235.29 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 152.135 236.06 152.505 ;
      VIA 235.29 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 146.715 236.08 147.045 ;
      VIA 235.29 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 146.695 236.06 147.065 ;
      VIA 235.29 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 141.275 236.08 141.605 ;
      VIA 235.29 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 141.255 236.06 141.625 ;
      VIA 235.29 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 135.835 236.08 136.165 ;
      VIA 235.29 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 135.815 236.06 136.185 ;
      VIA 235.29 136 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 130.395 236.08 130.725 ;
      VIA 235.29 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 130.375 236.06 130.745 ;
      VIA 235.29 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 124.955 236.08 125.285 ;
      VIA 235.29 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 124.935 236.06 125.305 ;
      VIA 235.29 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 119.515 236.08 119.845 ;
      VIA 235.29 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 119.495 236.06 119.865 ;
      VIA 235.29 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 114.075 236.08 114.405 ;
      VIA 235.29 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 114.055 236.06 114.425 ;
      VIA 235.29 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 108.635 236.08 108.965 ;
      VIA 235.29 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 108.615 236.06 108.985 ;
      VIA 235.29 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 103.195 236.08 103.525 ;
      VIA 235.29 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 103.175 236.06 103.545 ;
      VIA 235.29 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 97.755 236.08 98.085 ;
      VIA 235.29 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 97.735 236.06 98.105 ;
      VIA 235.29 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 92.315 236.08 92.645 ;
      VIA 235.29 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 92.295 236.06 92.665 ;
      VIA 235.29 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 86.875 236.08 87.205 ;
      VIA 235.29 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 86.855 236.06 87.225 ;
      VIA 235.29 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 81.435 236.08 81.765 ;
      VIA 235.29 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 81.415 236.06 81.785 ;
      VIA 235.29 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 75.995 236.08 76.325 ;
      VIA 235.29 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 75.975 236.06 76.345 ;
      VIA 235.29 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 70.555 236.08 70.885 ;
      VIA 235.29 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 70.535 236.06 70.905 ;
      VIA 235.29 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 65.115 236.08 65.445 ;
      VIA 235.29 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 65.095 236.06 65.465 ;
      VIA 235.29 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 59.675 236.08 60.005 ;
      VIA 235.29 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 59.655 236.06 60.025 ;
      VIA 235.29 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 54.235 236.08 54.565 ;
      VIA 235.29 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 54.215 236.06 54.585 ;
      VIA 235.29 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 48.795 236.08 49.125 ;
      VIA 235.29 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 48.775 236.06 49.145 ;
      VIA 235.29 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 43.355 236.08 43.685 ;
      VIA 235.29 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 43.335 236.06 43.705 ;
      VIA 235.29 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 37.915 236.08 38.245 ;
      VIA 235.29 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 37.895 236.06 38.265 ;
      VIA 235.29 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 32.475 236.08 32.805 ;
      VIA 235.29 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 32.455 236.06 32.825 ;
      VIA 235.29 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 27.035 236.08 27.365 ;
      VIA 235.29 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 27.015 236.06 27.385 ;
      VIA 235.29 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 21.595 236.08 21.925 ;
      VIA 235.29 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 21.575 236.06 21.945 ;
      VIA 235.29 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 16.155 236.08 16.485 ;
      VIA 235.29 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 16.135 236.06 16.505 ;
      VIA 235.29 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 10.715 236.08 11.045 ;
      VIA 235.29 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 10.695 236.06 11.065 ;
      VIA 235.29 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  234.5 5.275 236.08 5.605 ;
      VIA 235.29 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  234.52 5.255 236.06 5.625 ;
      VIA 235.29 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 235.29 5.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 282.715 208.94 283.045 ;
      VIA 208.15 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 282.695 208.92 283.065 ;
      VIA 208.15 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 277.275 208.94 277.605 ;
      VIA 208.15 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 277.255 208.92 277.625 ;
      VIA 208.15 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 271.835 208.94 272.165 ;
      VIA 208.15 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 271.815 208.92 272.185 ;
      VIA 208.15 272 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 266.395 208.94 266.725 ;
      VIA 208.15 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 266.375 208.92 266.745 ;
      VIA 208.15 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 260.955 208.94 261.285 ;
      VIA 208.15 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 260.935 208.92 261.305 ;
      VIA 208.15 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 255.515 208.94 255.845 ;
      VIA 208.15 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 255.495 208.92 255.865 ;
      VIA 208.15 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 250.075 208.94 250.405 ;
      VIA 208.15 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 250.055 208.92 250.425 ;
      VIA 208.15 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 244.635 208.94 244.965 ;
      VIA 208.15 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 244.615 208.92 244.985 ;
      VIA 208.15 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 239.195 208.94 239.525 ;
      VIA 208.15 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 239.175 208.92 239.545 ;
      VIA 208.15 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 233.755 208.94 234.085 ;
      VIA 208.15 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 233.735 208.92 234.105 ;
      VIA 208.15 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 228.315 208.94 228.645 ;
      VIA 208.15 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 228.295 208.92 228.665 ;
      VIA 208.15 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 222.875 208.94 223.205 ;
      VIA 208.15 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 222.855 208.92 223.225 ;
      VIA 208.15 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 217.435 208.94 217.765 ;
      VIA 208.15 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 217.415 208.92 217.785 ;
      VIA 208.15 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 211.995 208.94 212.325 ;
      VIA 208.15 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 211.975 208.92 212.345 ;
      VIA 208.15 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 206.555 208.94 206.885 ;
      VIA 208.15 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 206.535 208.92 206.905 ;
      VIA 208.15 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 201.115 208.94 201.445 ;
      VIA 208.15 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 201.095 208.92 201.465 ;
      VIA 208.15 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 195.675 208.94 196.005 ;
      VIA 208.15 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 195.655 208.92 196.025 ;
      VIA 208.15 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 190.235 208.94 190.565 ;
      VIA 208.15 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 190.215 208.92 190.585 ;
      VIA 208.15 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 184.795 208.94 185.125 ;
      VIA 208.15 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 184.775 208.92 185.145 ;
      VIA 208.15 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 179.355 208.94 179.685 ;
      VIA 208.15 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 179.335 208.92 179.705 ;
      VIA 208.15 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 173.915 208.94 174.245 ;
      VIA 208.15 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 173.895 208.92 174.265 ;
      VIA 208.15 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 168.475 208.94 168.805 ;
      VIA 208.15 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 168.455 208.92 168.825 ;
      VIA 208.15 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 163.035 208.94 163.365 ;
      VIA 208.15 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 163.015 208.92 163.385 ;
      VIA 208.15 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 157.595 208.94 157.925 ;
      VIA 208.15 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 157.575 208.92 157.945 ;
      VIA 208.15 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 152.155 208.94 152.485 ;
      VIA 208.15 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 152.135 208.92 152.505 ;
      VIA 208.15 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 146.715 208.94 147.045 ;
      VIA 208.15 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 146.695 208.92 147.065 ;
      VIA 208.15 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 141.275 208.94 141.605 ;
      VIA 208.15 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 141.255 208.92 141.625 ;
      VIA 208.15 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 135.835 208.94 136.165 ;
      VIA 208.15 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 135.815 208.92 136.185 ;
      VIA 208.15 136 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 130.395 208.94 130.725 ;
      VIA 208.15 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 130.375 208.92 130.745 ;
      VIA 208.15 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 124.955 208.94 125.285 ;
      VIA 208.15 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 124.935 208.92 125.305 ;
      VIA 208.15 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 119.515 208.94 119.845 ;
      VIA 208.15 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 119.495 208.92 119.865 ;
      VIA 208.15 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 114.075 208.94 114.405 ;
      VIA 208.15 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 114.055 208.92 114.425 ;
      VIA 208.15 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 108.635 208.94 108.965 ;
      VIA 208.15 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 108.615 208.92 108.985 ;
      VIA 208.15 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 103.195 208.94 103.525 ;
      VIA 208.15 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 103.175 208.92 103.545 ;
      VIA 208.15 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 97.755 208.94 98.085 ;
      VIA 208.15 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 97.735 208.92 98.105 ;
      VIA 208.15 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 92.315 208.94 92.645 ;
      VIA 208.15 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 92.295 208.92 92.665 ;
      VIA 208.15 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 86.875 208.94 87.205 ;
      VIA 208.15 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 86.855 208.92 87.225 ;
      VIA 208.15 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 81.435 208.94 81.765 ;
      VIA 208.15 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 81.415 208.92 81.785 ;
      VIA 208.15 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 75.995 208.94 76.325 ;
      VIA 208.15 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 75.975 208.92 76.345 ;
      VIA 208.15 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 70.555 208.94 70.885 ;
      VIA 208.15 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 70.535 208.92 70.905 ;
      VIA 208.15 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 65.115 208.94 65.445 ;
      VIA 208.15 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 65.095 208.92 65.465 ;
      VIA 208.15 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 59.675 208.94 60.005 ;
      VIA 208.15 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 59.655 208.92 60.025 ;
      VIA 208.15 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 54.235 208.94 54.565 ;
      VIA 208.15 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 54.215 208.92 54.585 ;
      VIA 208.15 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 48.795 208.94 49.125 ;
      VIA 208.15 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 48.775 208.92 49.145 ;
      VIA 208.15 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 43.355 208.94 43.685 ;
      VIA 208.15 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 43.335 208.92 43.705 ;
      VIA 208.15 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 37.915 208.94 38.245 ;
      VIA 208.15 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 37.895 208.92 38.265 ;
      VIA 208.15 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 32.475 208.94 32.805 ;
      VIA 208.15 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 32.455 208.92 32.825 ;
      VIA 208.15 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 27.035 208.94 27.365 ;
      VIA 208.15 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 27.015 208.92 27.385 ;
      VIA 208.15 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 21.595 208.94 21.925 ;
      VIA 208.15 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 21.575 208.92 21.945 ;
      VIA 208.15 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 16.155 208.94 16.485 ;
      VIA 208.15 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 16.135 208.92 16.505 ;
      VIA 208.15 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 10.715 208.94 11.045 ;
      VIA 208.15 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 10.695 208.92 11.065 ;
      VIA 208.15 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  207.36 5.275 208.94 5.605 ;
      VIA 208.15 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  207.38 5.255 208.92 5.625 ;
      VIA 208.15 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 208.15 5.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 282.715 181.8 283.045 ;
      VIA 181.01 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 282.695 181.78 283.065 ;
      VIA 181.01 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 277.275 181.8 277.605 ;
      VIA 181.01 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 277.255 181.78 277.625 ;
      VIA 181.01 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 271.835 181.8 272.165 ;
      VIA 181.01 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 271.815 181.78 272.185 ;
      VIA 181.01 272 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 266.395 181.8 266.725 ;
      VIA 181.01 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 266.375 181.78 266.745 ;
      VIA 181.01 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 260.955 181.8 261.285 ;
      VIA 181.01 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 260.935 181.78 261.305 ;
      VIA 181.01 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 255.515 181.8 255.845 ;
      VIA 181.01 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 255.495 181.78 255.865 ;
      VIA 181.01 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 250.075 181.8 250.405 ;
      VIA 181.01 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 250.055 181.78 250.425 ;
      VIA 181.01 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 244.635 181.8 244.965 ;
      VIA 181.01 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 244.615 181.78 244.985 ;
      VIA 181.01 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 239.195 181.8 239.525 ;
      VIA 181.01 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 239.175 181.78 239.545 ;
      VIA 181.01 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 233.755 181.8 234.085 ;
      VIA 181.01 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 233.735 181.78 234.105 ;
      VIA 181.01 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 228.315 181.8 228.645 ;
      VIA 181.01 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 228.295 181.78 228.665 ;
      VIA 181.01 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 222.875 181.8 223.205 ;
      VIA 181.01 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 222.855 181.78 223.225 ;
      VIA 181.01 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 217.435 181.8 217.765 ;
      VIA 181.01 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 217.415 181.78 217.785 ;
      VIA 181.01 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 211.995 181.8 212.325 ;
      VIA 181.01 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 211.975 181.78 212.345 ;
      VIA 181.01 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 206.555 181.8 206.885 ;
      VIA 181.01 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 206.535 181.78 206.905 ;
      VIA 181.01 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 201.115 181.8 201.445 ;
      VIA 181.01 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 201.095 181.78 201.465 ;
      VIA 181.01 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 195.675 181.8 196.005 ;
      VIA 181.01 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 195.655 181.78 196.025 ;
      VIA 181.01 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 190.235 181.8 190.565 ;
      VIA 181.01 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 190.215 181.78 190.585 ;
      VIA 181.01 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 184.795 181.8 185.125 ;
      VIA 181.01 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 184.775 181.78 185.145 ;
      VIA 181.01 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 179.355 181.8 179.685 ;
      VIA 181.01 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 179.335 181.78 179.705 ;
      VIA 181.01 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 173.915 181.8 174.245 ;
      VIA 181.01 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 173.895 181.78 174.265 ;
      VIA 181.01 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 168.475 181.8 168.805 ;
      VIA 181.01 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 168.455 181.78 168.825 ;
      VIA 181.01 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 163.035 181.8 163.365 ;
      VIA 181.01 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 163.015 181.78 163.385 ;
      VIA 181.01 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 157.595 181.8 157.925 ;
      VIA 181.01 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 157.575 181.78 157.945 ;
      VIA 181.01 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 152.155 181.8 152.485 ;
      VIA 181.01 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 152.135 181.78 152.505 ;
      VIA 181.01 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 146.715 181.8 147.045 ;
      VIA 181.01 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 146.695 181.78 147.065 ;
      VIA 181.01 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 141.275 181.8 141.605 ;
      VIA 181.01 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 141.255 181.78 141.625 ;
      VIA 181.01 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 135.835 181.8 136.165 ;
      VIA 181.01 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 135.815 181.78 136.185 ;
      VIA 181.01 136 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 130.395 181.8 130.725 ;
      VIA 181.01 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 130.375 181.78 130.745 ;
      VIA 181.01 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 124.955 181.8 125.285 ;
      VIA 181.01 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 124.935 181.78 125.305 ;
      VIA 181.01 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 119.515 181.8 119.845 ;
      VIA 181.01 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 119.495 181.78 119.865 ;
      VIA 181.01 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 114.075 181.8 114.405 ;
      VIA 181.01 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 114.055 181.78 114.425 ;
      VIA 181.01 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 108.635 181.8 108.965 ;
      VIA 181.01 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 108.615 181.78 108.985 ;
      VIA 181.01 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 103.195 181.8 103.525 ;
      VIA 181.01 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 103.175 181.78 103.545 ;
      VIA 181.01 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 97.755 181.8 98.085 ;
      VIA 181.01 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 97.735 181.78 98.105 ;
      VIA 181.01 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 92.315 181.8 92.645 ;
      VIA 181.01 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 92.295 181.78 92.665 ;
      VIA 181.01 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 86.875 181.8 87.205 ;
      VIA 181.01 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 86.855 181.78 87.225 ;
      VIA 181.01 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 81.435 181.8 81.765 ;
      VIA 181.01 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 81.415 181.78 81.785 ;
      VIA 181.01 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 75.995 181.8 76.325 ;
      VIA 181.01 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 75.975 181.78 76.345 ;
      VIA 181.01 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 70.555 181.8 70.885 ;
      VIA 181.01 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 70.535 181.78 70.905 ;
      VIA 181.01 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 65.115 181.8 65.445 ;
      VIA 181.01 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 65.095 181.78 65.465 ;
      VIA 181.01 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 59.675 181.8 60.005 ;
      VIA 181.01 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 59.655 181.78 60.025 ;
      VIA 181.01 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 54.235 181.8 54.565 ;
      VIA 181.01 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 54.215 181.78 54.585 ;
      VIA 181.01 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 48.795 181.8 49.125 ;
      VIA 181.01 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 48.775 181.78 49.145 ;
      VIA 181.01 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 43.355 181.8 43.685 ;
      VIA 181.01 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 43.335 181.78 43.705 ;
      VIA 181.01 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 37.915 181.8 38.245 ;
      VIA 181.01 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 37.895 181.78 38.265 ;
      VIA 181.01 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 32.475 181.8 32.805 ;
      VIA 181.01 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 32.455 181.78 32.825 ;
      VIA 181.01 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 27.035 181.8 27.365 ;
      VIA 181.01 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 27.015 181.78 27.385 ;
      VIA 181.01 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 21.595 181.8 21.925 ;
      VIA 181.01 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 21.575 181.78 21.945 ;
      VIA 181.01 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 16.155 181.8 16.485 ;
      VIA 181.01 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 16.135 181.78 16.505 ;
      VIA 181.01 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 10.715 181.8 11.045 ;
      VIA 181.01 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 10.695 181.78 11.065 ;
      VIA 181.01 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  180.22 5.275 181.8 5.605 ;
      VIA 181.01 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  180.24 5.255 181.78 5.625 ;
      VIA 181.01 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 181.01 5.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 282.715 154.66 283.045 ;
      VIA 153.87 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 282.695 154.64 283.065 ;
      VIA 153.87 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 277.275 154.66 277.605 ;
      VIA 153.87 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 277.255 154.64 277.625 ;
      VIA 153.87 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 271.835 154.66 272.165 ;
      VIA 153.87 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 271.815 154.64 272.185 ;
      VIA 153.87 272 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 266.395 154.66 266.725 ;
      VIA 153.87 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 266.375 154.64 266.745 ;
      VIA 153.87 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 260.955 154.66 261.285 ;
      VIA 153.87 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 260.935 154.64 261.305 ;
      VIA 153.87 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 255.515 154.66 255.845 ;
      VIA 153.87 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 255.495 154.64 255.865 ;
      VIA 153.87 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 250.075 154.66 250.405 ;
      VIA 153.87 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 250.055 154.64 250.425 ;
      VIA 153.87 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 244.635 154.66 244.965 ;
      VIA 153.87 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 244.615 154.64 244.985 ;
      VIA 153.87 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 239.195 154.66 239.525 ;
      VIA 153.87 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 239.175 154.64 239.545 ;
      VIA 153.87 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 233.755 154.66 234.085 ;
      VIA 153.87 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 233.735 154.64 234.105 ;
      VIA 153.87 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 228.315 154.66 228.645 ;
      VIA 153.87 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 228.295 154.64 228.665 ;
      VIA 153.87 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 222.875 154.66 223.205 ;
      VIA 153.87 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 222.855 154.64 223.225 ;
      VIA 153.87 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 217.435 154.66 217.765 ;
      VIA 153.87 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 217.415 154.64 217.785 ;
      VIA 153.87 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 211.995 154.66 212.325 ;
      VIA 153.87 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 211.975 154.64 212.345 ;
      VIA 153.87 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 206.555 154.66 206.885 ;
      VIA 153.87 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 206.535 154.64 206.905 ;
      VIA 153.87 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 201.115 154.66 201.445 ;
      VIA 153.87 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 201.095 154.64 201.465 ;
      VIA 153.87 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 195.675 154.66 196.005 ;
      VIA 153.87 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 195.655 154.64 196.025 ;
      VIA 153.87 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 190.235 154.66 190.565 ;
      VIA 153.87 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 190.215 154.64 190.585 ;
      VIA 153.87 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 184.795 154.66 185.125 ;
      VIA 153.87 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 184.775 154.64 185.145 ;
      VIA 153.87 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 179.355 154.66 179.685 ;
      VIA 153.87 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 179.335 154.64 179.705 ;
      VIA 153.87 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 173.915 154.66 174.245 ;
      VIA 153.87 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 173.895 154.64 174.265 ;
      VIA 153.87 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 168.475 154.66 168.805 ;
      VIA 153.87 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 168.455 154.64 168.825 ;
      VIA 153.87 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 163.035 154.66 163.365 ;
      VIA 153.87 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 163.015 154.64 163.385 ;
      VIA 153.87 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 157.595 154.66 157.925 ;
      VIA 153.87 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 157.575 154.64 157.945 ;
      VIA 153.87 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 152.155 154.66 152.485 ;
      VIA 153.87 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 152.135 154.64 152.505 ;
      VIA 153.87 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 146.715 154.66 147.045 ;
      VIA 153.87 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 146.695 154.64 147.065 ;
      VIA 153.87 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 141.275 154.66 141.605 ;
      VIA 153.87 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 141.255 154.64 141.625 ;
      VIA 153.87 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 135.835 154.66 136.165 ;
      VIA 153.87 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 135.815 154.64 136.185 ;
      VIA 153.87 136 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 130.395 154.66 130.725 ;
      VIA 153.87 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 130.375 154.64 130.745 ;
      VIA 153.87 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 124.955 154.66 125.285 ;
      VIA 153.87 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 124.935 154.64 125.305 ;
      VIA 153.87 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 119.515 154.66 119.845 ;
      VIA 153.87 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 119.495 154.64 119.865 ;
      VIA 153.87 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 114.075 154.66 114.405 ;
      VIA 153.87 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 114.055 154.64 114.425 ;
      VIA 153.87 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 108.635 154.66 108.965 ;
      VIA 153.87 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 108.615 154.64 108.985 ;
      VIA 153.87 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 103.195 154.66 103.525 ;
      VIA 153.87 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 103.175 154.64 103.545 ;
      VIA 153.87 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 97.755 154.66 98.085 ;
      VIA 153.87 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 97.735 154.64 98.105 ;
      VIA 153.87 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 92.315 154.66 92.645 ;
      VIA 153.87 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 92.295 154.64 92.665 ;
      VIA 153.87 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 86.875 154.66 87.205 ;
      VIA 153.87 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 86.855 154.64 87.225 ;
      VIA 153.87 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 81.435 154.66 81.765 ;
      VIA 153.87 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 81.415 154.64 81.785 ;
      VIA 153.87 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 75.995 154.66 76.325 ;
      VIA 153.87 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 75.975 154.64 76.345 ;
      VIA 153.87 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 70.555 154.66 70.885 ;
      VIA 153.87 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 70.535 154.64 70.905 ;
      VIA 153.87 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 65.115 154.66 65.445 ;
      VIA 153.87 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 65.095 154.64 65.465 ;
      VIA 153.87 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 59.675 154.66 60.005 ;
      VIA 153.87 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 59.655 154.64 60.025 ;
      VIA 153.87 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 54.235 154.66 54.565 ;
      VIA 153.87 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 54.215 154.64 54.585 ;
      VIA 153.87 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 48.795 154.66 49.125 ;
      VIA 153.87 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 48.775 154.64 49.145 ;
      VIA 153.87 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 43.355 154.66 43.685 ;
      VIA 153.87 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 43.335 154.64 43.705 ;
      VIA 153.87 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 37.915 154.66 38.245 ;
      VIA 153.87 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 37.895 154.64 38.265 ;
      VIA 153.87 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 32.475 154.66 32.805 ;
      VIA 153.87 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 32.455 154.64 32.825 ;
      VIA 153.87 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 27.035 154.66 27.365 ;
      VIA 153.87 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 27.015 154.64 27.385 ;
      VIA 153.87 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 21.595 154.66 21.925 ;
      VIA 153.87 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 21.575 154.64 21.945 ;
      VIA 153.87 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 16.155 154.66 16.485 ;
      VIA 153.87 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 16.135 154.64 16.505 ;
      VIA 153.87 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 10.715 154.66 11.045 ;
      VIA 153.87 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 10.695 154.64 11.065 ;
      VIA 153.87 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  153.08 5.275 154.66 5.605 ;
      VIA 153.87 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  153.1 5.255 154.64 5.625 ;
      VIA 153.87 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 153.87 5.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 282.715 127.52 283.045 ;
      VIA 126.73 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 282.695 127.5 283.065 ;
      VIA 126.73 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 277.275 127.52 277.605 ;
      VIA 126.73 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 277.255 127.5 277.625 ;
      VIA 126.73 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 271.835 127.52 272.165 ;
      VIA 126.73 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 271.815 127.5 272.185 ;
      VIA 126.73 272 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 266.395 127.52 266.725 ;
      VIA 126.73 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 266.375 127.5 266.745 ;
      VIA 126.73 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 260.955 127.52 261.285 ;
      VIA 126.73 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 260.935 127.5 261.305 ;
      VIA 126.73 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 255.515 127.52 255.845 ;
      VIA 126.73 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 255.495 127.5 255.865 ;
      VIA 126.73 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 250.075 127.52 250.405 ;
      VIA 126.73 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 250.055 127.5 250.425 ;
      VIA 126.73 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 244.635 127.52 244.965 ;
      VIA 126.73 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 244.615 127.5 244.985 ;
      VIA 126.73 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 239.195 127.52 239.525 ;
      VIA 126.73 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 239.175 127.5 239.545 ;
      VIA 126.73 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 233.755 127.52 234.085 ;
      VIA 126.73 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 233.735 127.5 234.105 ;
      VIA 126.73 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 228.315 127.52 228.645 ;
      VIA 126.73 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 228.295 127.5 228.665 ;
      VIA 126.73 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 222.875 127.52 223.205 ;
      VIA 126.73 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 222.855 127.5 223.225 ;
      VIA 126.73 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 217.435 127.52 217.765 ;
      VIA 126.73 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 217.415 127.5 217.785 ;
      VIA 126.73 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 211.995 127.52 212.325 ;
      VIA 126.73 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 211.975 127.5 212.345 ;
      VIA 126.73 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 206.555 127.52 206.885 ;
      VIA 126.73 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 206.535 127.5 206.905 ;
      VIA 126.73 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 201.115 127.52 201.445 ;
      VIA 126.73 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 201.095 127.5 201.465 ;
      VIA 126.73 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 195.675 127.52 196.005 ;
      VIA 126.73 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 195.655 127.5 196.025 ;
      VIA 126.73 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 190.235 127.52 190.565 ;
      VIA 126.73 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 190.215 127.5 190.585 ;
      VIA 126.73 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 184.795 127.52 185.125 ;
      VIA 126.73 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 184.775 127.5 185.145 ;
      VIA 126.73 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 179.355 127.52 179.685 ;
      VIA 126.73 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 179.335 127.5 179.705 ;
      VIA 126.73 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 173.915 127.52 174.245 ;
      VIA 126.73 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 173.895 127.5 174.265 ;
      VIA 126.73 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 168.475 127.52 168.805 ;
      VIA 126.73 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 168.455 127.5 168.825 ;
      VIA 126.73 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 163.035 127.52 163.365 ;
      VIA 126.73 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 163.015 127.5 163.385 ;
      VIA 126.73 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 157.595 127.52 157.925 ;
      VIA 126.73 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 157.575 127.5 157.945 ;
      VIA 126.73 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 152.155 127.52 152.485 ;
      VIA 126.73 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 152.135 127.5 152.505 ;
      VIA 126.73 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 146.715 127.52 147.045 ;
      VIA 126.73 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 146.695 127.5 147.065 ;
      VIA 126.73 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 141.275 127.52 141.605 ;
      VIA 126.73 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 141.255 127.5 141.625 ;
      VIA 126.73 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 135.835 127.52 136.165 ;
      VIA 126.73 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 135.815 127.5 136.185 ;
      VIA 126.73 136 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 130.395 127.52 130.725 ;
      VIA 126.73 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 130.375 127.5 130.745 ;
      VIA 126.73 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 124.955 127.52 125.285 ;
      VIA 126.73 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 124.935 127.5 125.305 ;
      VIA 126.73 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 119.515 127.52 119.845 ;
      VIA 126.73 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 119.495 127.5 119.865 ;
      VIA 126.73 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 114.075 127.52 114.405 ;
      VIA 126.73 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 114.055 127.5 114.425 ;
      VIA 126.73 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 108.635 127.52 108.965 ;
      VIA 126.73 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 108.615 127.5 108.985 ;
      VIA 126.73 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 103.195 127.52 103.525 ;
      VIA 126.73 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 103.175 127.5 103.545 ;
      VIA 126.73 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 97.755 127.52 98.085 ;
      VIA 126.73 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 97.735 127.5 98.105 ;
      VIA 126.73 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 92.315 127.52 92.645 ;
      VIA 126.73 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 92.295 127.5 92.665 ;
      VIA 126.73 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 86.875 127.52 87.205 ;
      VIA 126.73 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 86.855 127.5 87.225 ;
      VIA 126.73 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 81.435 127.52 81.765 ;
      VIA 126.73 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 81.415 127.5 81.785 ;
      VIA 126.73 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 75.995 127.52 76.325 ;
      VIA 126.73 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 75.975 127.5 76.345 ;
      VIA 126.73 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 70.555 127.52 70.885 ;
      VIA 126.73 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 70.535 127.5 70.905 ;
      VIA 126.73 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 65.115 127.52 65.445 ;
      VIA 126.73 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 65.095 127.5 65.465 ;
      VIA 126.73 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 59.675 127.52 60.005 ;
      VIA 126.73 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 59.655 127.5 60.025 ;
      VIA 126.73 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 54.235 127.52 54.565 ;
      VIA 126.73 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 54.215 127.5 54.585 ;
      VIA 126.73 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 48.795 127.52 49.125 ;
      VIA 126.73 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 48.775 127.5 49.145 ;
      VIA 126.73 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 43.355 127.52 43.685 ;
      VIA 126.73 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 43.335 127.5 43.705 ;
      VIA 126.73 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 37.915 127.52 38.245 ;
      VIA 126.73 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 37.895 127.5 38.265 ;
      VIA 126.73 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 32.475 127.52 32.805 ;
      VIA 126.73 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 32.455 127.5 32.825 ;
      VIA 126.73 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 27.035 127.52 27.365 ;
      VIA 126.73 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 27.015 127.5 27.385 ;
      VIA 126.73 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 21.595 127.52 21.925 ;
      VIA 126.73 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 21.575 127.5 21.945 ;
      VIA 126.73 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 16.155 127.52 16.485 ;
      VIA 126.73 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 16.135 127.5 16.505 ;
      VIA 126.73 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 10.715 127.52 11.045 ;
      VIA 126.73 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 10.695 127.5 11.065 ;
      VIA 126.73 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  125.94 5.275 127.52 5.605 ;
      VIA 126.73 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  125.96 5.255 127.5 5.625 ;
      VIA 126.73 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 126.73 5.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 282.715 100.38 283.045 ;
      VIA 99.59 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 282.695 100.36 283.065 ;
      VIA 99.59 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 277.275 100.38 277.605 ;
      VIA 99.59 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 277.255 100.36 277.625 ;
      VIA 99.59 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 271.835 100.38 272.165 ;
      VIA 99.59 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 271.815 100.36 272.185 ;
      VIA 99.59 272 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 266.395 100.38 266.725 ;
      VIA 99.59 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 266.375 100.36 266.745 ;
      VIA 99.59 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 260.955 100.38 261.285 ;
      VIA 99.59 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 260.935 100.36 261.305 ;
      VIA 99.59 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 255.515 100.38 255.845 ;
      VIA 99.59 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 255.495 100.36 255.865 ;
      VIA 99.59 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 250.075 100.38 250.405 ;
      VIA 99.59 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 250.055 100.36 250.425 ;
      VIA 99.59 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 244.635 100.38 244.965 ;
      VIA 99.59 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 244.615 100.36 244.985 ;
      VIA 99.59 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 239.195 100.38 239.525 ;
      VIA 99.59 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 239.175 100.36 239.545 ;
      VIA 99.59 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 233.755 100.38 234.085 ;
      VIA 99.59 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 233.735 100.36 234.105 ;
      VIA 99.59 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 228.315 100.38 228.645 ;
      VIA 99.59 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 228.295 100.36 228.665 ;
      VIA 99.59 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 222.875 100.38 223.205 ;
      VIA 99.59 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 222.855 100.36 223.225 ;
      VIA 99.59 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 217.435 100.38 217.765 ;
      VIA 99.59 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 217.415 100.36 217.785 ;
      VIA 99.59 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 211.995 100.38 212.325 ;
      VIA 99.59 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 211.975 100.36 212.345 ;
      VIA 99.59 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 206.555 100.38 206.885 ;
      VIA 99.59 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 206.535 100.36 206.905 ;
      VIA 99.59 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 201.115 100.38 201.445 ;
      VIA 99.59 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 201.095 100.36 201.465 ;
      VIA 99.59 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 195.675 100.38 196.005 ;
      VIA 99.59 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 195.655 100.36 196.025 ;
      VIA 99.59 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 190.235 100.38 190.565 ;
      VIA 99.59 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 190.215 100.36 190.585 ;
      VIA 99.59 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 184.795 100.38 185.125 ;
      VIA 99.59 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 184.775 100.36 185.145 ;
      VIA 99.59 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 179.355 100.38 179.685 ;
      VIA 99.59 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 179.335 100.36 179.705 ;
      VIA 99.59 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 173.915 100.38 174.245 ;
      VIA 99.59 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 173.895 100.36 174.265 ;
      VIA 99.59 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 168.475 100.38 168.805 ;
      VIA 99.59 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 168.455 100.36 168.825 ;
      VIA 99.59 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 163.035 100.38 163.365 ;
      VIA 99.59 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 163.015 100.36 163.385 ;
      VIA 99.59 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 157.595 100.38 157.925 ;
      VIA 99.59 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 157.575 100.36 157.945 ;
      VIA 99.59 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 152.155 100.38 152.485 ;
      VIA 99.59 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 152.135 100.36 152.505 ;
      VIA 99.59 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 146.715 100.38 147.045 ;
      VIA 99.59 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 146.695 100.36 147.065 ;
      VIA 99.59 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 141.275 100.38 141.605 ;
      VIA 99.59 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 141.255 100.36 141.625 ;
      VIA 99.59 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 135.835 100.38 136.165 ;
      VIA 99.59 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 135.815 100.36 136.185 ;
      VIA 99.59 136 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 130.395 100.38 130.725 ;
      VIA 99.59 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 130.375 100.36 130.745 ;
      VIA 99.59 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 124.955 100.38 125.285 ;
      VIA 99.59 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 124.935 100.36 125.305 ;
      VIA 99.59 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 119.515 100.38 119.845 ;
      VIA 99.59 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 119.495 100.36 119.865 ;
      VIA 99.59 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 114.075 100.38 114.405 ;
      VIA 99.59 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 114.055 100.36 114.425 ;
      VIA 99.59 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 108.635 100.38 108.965 ;
      VIA 99.59 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 108.615 100.36 108.985 ;
      VIA 99.59 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 103.195 100.38 103.525 ;
      VIA 99.59 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 103.175 100.36 103.545 ;
      VIA 99.59 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 97.755 100.38 98.085 ;
      VIA 99.59 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 97.735 100.36 98.105 ;
      VIA 99.59 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 92.315 100.38 92.645 ;
      VIA 99.59 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 92.295 100.36 92.665 ;
      VIA 99.59 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 86.875 100.38 87.205 ;
      VIA 99.59 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 86.855 100.36 87.225 ;
      VIA 99.59 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 81.435 100.38 81.765 ;
      VIA 99.59 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 81.415 100.36 81.785 ;
      VIA 99.59 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 75.995 100.38 76.325 ;
      VIA 99.59 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 75.975 100.36 76.345 ;
      VIA 99.59 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 70.555 100.38 70.885 ;
      VIA 99.59 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 70.535 100.36 70.905 ;
      VIA 99.59 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 65.115 100.38 65.445 ;
      VIA 99.59 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 65.095 100.36 65.465 ;
      VIA 99.59 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 59.675 100.38 60.005 ;
      VIA 99.59 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 59.655 100.36 60.025 ;
      VIA 99.59 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 54.235 100.38 54.565 ;
      VIA 99.59 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 54.215 100.36 54.585 ;
      VIA 99.59 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 48.795 100.38 49.125 ;
      VIA 99.59 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 48.775 100.36 49.145 ;
      VIA 99.59 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 43.355 100.38 43.685 ;
      VIA 99.59 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 43.335 100.36 43.705 ;
      VIA 99.59 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 37.915 100.38 38.245 ;
      VIA 99.59 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 37.895 100.36 38.265 ;
      VIA 99.59 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 32.475 100.38 32.805 ;
      VIA 99.59 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 32.455 100.36 32.825 ;
      VIA 99.59 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 27.035 100.38 27.365 ;
      VIA 99.59 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 27.015 100.36 27.385 ;
      VIA 99.59 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 21.595 100.38 21.925 ;
      VIA 99.59 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 21.575 100.36 21.945 ;
      VIA 99.59 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 16.155 100.38 16.485 ;
      VIA 99.59 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 16.135 100.36 16.505 ;
      VIA 99.59 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 10.715 100.38 11.045 ;
      VIA 99.59 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 10.695 100.36 11.065 ;
      VIA 99.59 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  98.8 5.275 100.38 5.605 ;
      VIA 99.59 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  98.82 5.255 100.36 5.625 ;
      VIA 99.59 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 99.59 5.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 282.715 73.24 283.045 ;
      VIA 72.45 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 282.695 73.22 283.065 ;
      VIA 72.45 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 277.275 73.24 277.605 ;
      VIA 72.45 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 277.255 73.22 277.625 ;
      VIA 72.45 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 271.835 73.24 272.165 ;
      VIA 72.45 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 271.815 73.22 272.185 ;
      VIA 72.45 272 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 266.395 73.24 266.725 ;
      VIA 72.45 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 266.375 73.22 266.745 ;
      VIA 72.45 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 260.955 73.24 261.285 ;
      VIA 72.45 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 260.935 73.22 261.305 ;
      VIA 72.45 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 255.515 73.24 255.845 ;
      VIA 72.45 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 255.495 73.22 255.865 ;
      VIA 72.45 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 250.075 73.24 250.405 ;
      VIA 72.45 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 250.055 73.22 250.425 ;
      VIA 72.45 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 244.635 73.24 244.965 ;
      VIA 72.45 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 244.615 73.22 244.985 ;
      VIA 72.45 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 239.195 73.24 239.525 ;
      VIA 72.45 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 239.175 73.22 239.545 ;
      VIA 72.45 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 233.755 73.24 234.085 ;
      VIA 72.45 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 233.735 73.22 234.105 ;
      VIA 72.45 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 228.315 73.24 228.645 ;
      VIA 72.45 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 228.295 73.22 228.665 ;
      VIA 72.45 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 222.875 73.24 223.205 ;
      VIA 72.45 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 222.855 73.22 223.225 ;
      VIA 72.45 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 217.435 73.24 217.765 ;
      VIA 72.45 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 217.415 73.22 217.785 ;
      VIA 72.45 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 211.995 73.24 212.325 ;
      VIA 72.45 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 211.975 73.22 212.345 ;
      VIA 72.45 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 206.555 73.24 206.885 ;
      VIA 72.45 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 206.535 73.22 206.905 ;
      VIA 72.45 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 201.115 73.24 201.445 ;
      VIA 72.45 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 201.095 73.22 201.465 ;
      VIA 72.45 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 195.675 73.24 196.005 ;
      VIA 72.45 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 195.655 73.22 196.025 ;
      VIA 72.45 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 190.235 73.24 190.565 ;
      VIA 72.45 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 190.215 73.22 190.585 ;
      VIA 72.45 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 184.795 73.24 185.125 ;
      VIA 72.45 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 184.775 73.22 185.145 ;
      VIA 72.45 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 179.355 73.24 179.685 ;
      VIA 72.45 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 179.335 73.22 179.705 ;
      VIA 72.45 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 173.915 73.24 174.245 ;
      VIA 72.45 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 173.895 73.22 174.265 ;
      VIA 72.45 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 168.475 73.24 168.805 ;
      VIA 72.45 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 168.455 73.22 168.825 ;
      VIA 72.45 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 163.035 73.24 163.365 ;
      VIA 72.45 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 163.015 73.22 163.385 ;
      VIA 72.45 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 157.595 73.24 157.925 ;
      VIA 72.45 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 157.575 73.22 157.945 ;
      VIA 72.45 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 152.155 73.24 152.485 ;
      VIA 72.45 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 152.135 73.22 152.505 ;
      VIA 72.45 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 146.715 73.24 147.045 ;
      VIA 72.45 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 146.695 73.22 147.065 ;
      VIA 72.45 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 141.275 73.24 141.605 ;
      VIA 72.45 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 141.255 73.22 141.625 ;
      VIA 72.45 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 135.835 73.24 136.165 ;
      VIA 72.45 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 135.815 73.22 136.185 ;
      VIA 72.45 136 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 130.395 73.24 130.725 ;
      VIA 72.45 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 130.375 73.22 130.745 ;
      VIA 72.45 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 124.955 73.24 125.285 ;
      VIA 72.45 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 124.935 73.22 125.305 ;
      VIA 72.45 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 119.515 73.24 119.845 ;
      VIA 72.45 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 119.495 73.22 119.865 ;
      VIA 72.45 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 114.075 73.24 114.405 ;
      VIA 72.45 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 114.055 73.22 114.425 ;
      VIA 72.45 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 108.635 73.24 108.965 ;
      VIA 72.45 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 108.615 73.22 108.985 ;
      VIA 72.45 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 103.195 73.24 103.525 ;
      VIA 72.45 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 103.175 73.22 103.545 ;
      VIA 72.45 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 97.755 73.24 98.085 ;
      VIA 72.45 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 97.735 73.22 98.105 ;
      VIA 72.45 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 92.315 73.24 92.645 ;
      VIA 72.45 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 92.295 73.22 92.665 ;
      VIA 72.45 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 86.875 73.24 87.205 ;
      VIA 72.45 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 86.855 73.22 87.225 ;
      VIA 72.45 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 81.435 73.24 81.765 ;
      VIA 72.45 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 81.415 73.22 81.785 ;
      VIA 72.45 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 75.995 73.24 76.325 ;
      VIA 72.45 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 75.975 73.22 76.345 ;
      VIA 72.45 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 70.555 73.24 70.885 ;
      VIA 72.45 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 70.535 73.22 70.905 ;
      VIA 72.45 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 65.115 73.24 65.445 ;
      VIA 72.45 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 65.095 73.22 65.465 ;
      VIA 72.45 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 59.675 73.24 60.005 ;
      VIA 72.45 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 59.655 73.22 60.025 ;
      VIA 72.45 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 54.235 73.24 54.565 ;
      VIA 72.45 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 54.215 73.22 54.585 ;
      VIA 72.45 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 48.795 73.24 49.125 ;
      VIA 72.45 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 48.775 73.22 49.145 ;
      VIA 72.45 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 43.355 73.24 43.685 ;
      VIA 72.45 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 43.335 73.22 43.705 ;
      VIA 72.45 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 37.915 73.24 38.245 ;
      VIA 72.45 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 37.895 73.22 38.265 ;
      VIA 72.45 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 32.475 73.24 32.805 ;
      VIA 72.45 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 32.455 73.22 32.825 ;
      VIA 72.45 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 27.035 73.24 27.365 ;
      VIA 72.45 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 27.015 73.22 27.385 ;
      VIA 72.45 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 21.595 73.24 21.925 ;
      VIA 72.45 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 21.575 73.22 21.945 ;
      VIA 72.45 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 16.155 73.24 16.485 ;
      VIA 72.45 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 16.135 73.22 16.505 ;
      VIA 72.45 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 10.715 73.24 11.045 ;
      VIA 72.45 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 10.695 73.22 11.065 ;
      VIA 72.45 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  71.66 5.275 73.24 5.605 ;
      VIA 72.45 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  71.68 5.255 73.22 5.625 ;
      VIA 72.45 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 72.45 5.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 282.715 46.1 283.045 ;
      VIA 45.31 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 282.695 46.08 283.065 ;
      VIA 45.31 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 277.275 46.1 277.605 ;
      VIA 45.31 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 277.255 46.08 277.625 ;
      VIA 45.31 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 271.835 46.1 272.165 ;
      VIA 45.31 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 271.815 46.08 272.185 ;
      VIA 45.31 272 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 266.395 46.1 266.725 ;
      VIA 45.31 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 266.375 46.08 266.745 ;
      VIA 45.31 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 260.955 46.1 261.285 ;
      VIA 45.31 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 260.935 46.08 261.305 ;
      VIA 45.31 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 255.515 46.1 255.845 ;
      VIA 45.31 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 255.495 46.08 255.865 ;
      VIA 45.31 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 250.075 46.1 250.405 ;
      VIA 45.31 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 250.055 46.08 250.425 ;
      VIA 45.31 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 244.635 46.1 244.965 ;
      VIA 45.31 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 244.615 46.08 244.985 ;
      VIA 45.31 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 239.195 46.1 239.525 ;
      VIA 45.31 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 239.175 46.08 239.545 ;
      VIA 45.31 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 233.755 46.1 234.085 ;
      VIA 45.31 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 233.735 46.08 234.105 ;
      VIA 45.31 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 228.315 46.1 228.645 ;
      VIA 45.31 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 228.295 46.08 228.665 ;
      VIA 45.31 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 222.875 46.1 223.205 ;
      VIA 45.31 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 222.855 46.08 223.225 ;
      VIA 45.31 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 217.435 46.1 217.765 ;
      VIA 45.31 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 217.415 46.08 217.785 ;
      VIA 45.31 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 211.995 46.1 212.325 ;
      VIA 45.31 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 211.975 46.08 212.345 ;
      VIA 45.31 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 206.555 46.1 206.885 ;
      VIA 45.31 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 206.535 46.08 206.905 ;
      VIA 45.31 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 201.115 46.1 201.445 ;
      VIA 45.31 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 201.095 46.08 201.465 ;
      VIA 45.31 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 195.675 46.1 196.005 ;
      VIA 45.31 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 195.655 46.08 196.025 ;
      VIA 45.31 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 190.235 46.1 190.565 ;
      VIA 45.31 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 190.215 46.08 190.585 ;
      VIA 45.31 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 184.795 46.1 185.125 ;
      VIA 45.31 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 184.775 46.08 185.145 ;
      VIA 45.31 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 179.355 46.1 179.685 ;
      VIA 45.31 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 179.335 46.08 179.705 ;
      VIA 45.31 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 173.915 46.1 174.245 ;
      VIA 45.31 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 173.895 46.08 174.265 ;
      VIA 45.31 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 168.475 46.1 168.805 ;
      VIA 45.31 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 168.455 46.08 168.825 ;
      VIA 45.31 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 163.035 46.1 163.365 ;
      VIA 45.31 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 163.015 46.08 163.385 ;
      VIA 45.31 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 157.595 46.1 157.925 ;
      VIA 45.31 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 157.575 46.08 157.945 ;
      VIA 45.31 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 152.155 46.1 152.485 ;
      VIA 45.31 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 152.135 46.08 152.505 ;
      VIA 45.31 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 146.715 46.1 147.045 ;
      VIA 45.31 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 146.695 46.08 147.065 ;
      VIA 45.31 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 141.275 46.1 141.605 ;
      VIA 45.31 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 141.255 46.08 141.625 ;
      VIA 45.31 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 135.835 46.1 136.165 ;
      VIA 45.31 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 135.815 46.08 136.185 ;
      VIA 45.31 136 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 130.395 46.1 130.725 ;
      VIA 45.31 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 130.375 46.08 130.745 ;
      VIA 45.31 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 124.955 46.1 125.285 ;
      VIA 45.31 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 124.935 46.08 125.305 ;
      VIA 45.31 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 119.515 46.1 119.845 ;
      VIA 45.31 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 119.495 46.08 119.865 ;
      VIA 45.31 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 114.075 46.1 114.405 ;
      VIA 45.31 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 114.055 46.08 114.425 ;
      VIA 45.31 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 108.635 46.1 108.965 ;
      VIA 45.31 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 108.615 46.08 108.985 ;
      VIA 45.31 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 103.195 46.1 103.525 ;
      VIA 45.31 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 103.175 46.08 103.545 ;
      VIA 45.31 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 97.755 46.1 98.085 ;
      VIA 45.31 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 97.735 46.08 98.105 ;
      VIA 45.31 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 92.315 46.1 92.645 ;
      VIA 45.31 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 92.295 46.08 92.665 ;
      VIA 45.31 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 86.875 46.1 87.205 ;
      VIA 45.31 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 86.855 46.08 87.225 ;
      VIA 45.31 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 81.435 46.1 81.765 ;
      VIA 45.31 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 81.415 46.08 81.785 ;
      VIA 45.31 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 75.995 46.1 76.325 ;
      VIA 45.31 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 75.975 46.08 76.345 ;
      VIA 45.31 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 70.555 46.1 70.885 ;
      VIA 45.31 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 70.535 46.08 70.905 ;
      VIA 45.31 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 65.115 46.1 65.445 ;
      VIA 45.31 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 65.095 46.08 65.465 ;
      VIA 45.31 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 59.675 46.1 60.005 ;
      VIA 45.31 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 59.655 46.08 60.025 ;
      VIA 45.31 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 54.235 46.1 54.565 ;
      VIA 45.31 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 54.215 46.08 54.585 ;
      VIA 45.31 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 48.795 46.1 49.125 ;
      VIA 45.31 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 48.775 46.08 49.145 ;
      VIA 45.31 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 43.355 46.1 43.685 ;
      VIA 45.31 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 43.335 46.08 43.705 ;
      VIA 45.31 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 37.915 46.1 38.245 ;
      VIA 45.31 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 37.895 46.08 38.265 ;
      VIA 45.31 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 32.475 46.1 32.805 ;
      VIA 45.31 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 32.455 46.08 32.825 ;
      VIA 45.31 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 27.035 46.1 27.365 ;
      VIA 45.31 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 27.015 46.08 27.385 ;
      VIA 45.31 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 21.595 46.1 21.925 ;
      VIA 45.31 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 21.575 46.08 21.945 ;
      VIA 45.31 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 16.155 46.1 16.485 ;
      VIA 45.31 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 16.135 46.08 16.505 ;
      VIA 45.31 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 10.715 46.1 11.045 ;
      VIA 45.31 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 10.695 46.08 11.065 ;
      VIA 45.31 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  44.52 5.275 46.1 5.605 ;
      VIA 45.31 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  44.54 5.255 46.08 5.625 ;
      VIA 45.31 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 45.31 5.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 282.715 18.96 283.045 ;
      VIA 18.17 282.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 282.695 18.94 283.065 ;
      VIA 18.17 282.88 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 282.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 277.275 18.96 277.605 ;
      VIA 18.17 277.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 277.255 18.94 277.625 ;
      VIA 18.17 277.44 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 277.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 271.835 18.96 272.165 ;
      VIA 18.17 272 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 271.815 18.94 272.185 ;
      VIA 18.17 272 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 272 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 266.395 18.96 266.725 ;
      VIA 18.17 266.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 266.375 18.94 266.745 ;
      VIA 18.17 266.56 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 266.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 260.955 18.96 261.285 ;
      VIA 18.17 261.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 260.935 18.94 261.305 ;
      VIA 18.17 261.12 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 261.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 255.515 18.96 255.845 ;
      VIA 18.17 255.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 255.495 18.94 255.865 ;
      VIA 18.17 255.68 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 255.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 250.075 18.96 250.405 ;
      VIA 18.17 250.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 250.055 18.94 250.425 ;
      VIA 18.17 250.24 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 250.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 244.635 18.96 244.965 ;
      VIA 18.17 244.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 244.615 18.94 244.985 ;
      VIA 18.17 244.8 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 244.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 239.195 18.96 239.525 ;
      VIA 18.17 239.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 239.175 18.94 239.545 ;
      VIA 18.17 239.36 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 239.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 233.755 18.96 234.085 ;
      VIA 18.17 233.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 233.735 18.94 234.105 ;
      VIA 18.17 233.92 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 233.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 228.315 18.96 228.645 ;
      VIA 18.17 228.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 228.295 18.94 228.665 ;
      VIA 18.17 228.48 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 228.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 222.875 18.96 223.205 ;
      VIA 18.17 223.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 222.855 18.94 223.225 ;
      VIA 18.17 223.04 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 223.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 217.435 18.96 217.765 ;
      VIA 18.17 217.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 217.415 18.94 217.785 ;
      VIA 18.17 217.6 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 217.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 211.995 18.96 212.325 ;
      VIA 18.17 212.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 211.975 18.94 212.345 ;
      VIA 18.17 212.16 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 212.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 206.555 18.96 206.885 ;
      VIA 18.17 206.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 206.535 18.94 206.905 ;
      VIA 18.17 206.72 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 206.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 201.115 18.96 201.445 ;
      VIA 18.17 201.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 201.095 18.94 201.465 ;
      VIA 18.17 201.28 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 201.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 195.675 18.96 196.005 ;
      VIA 18.17 195.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 195.655 18.94 196.025 ;
      VIA 18.17 195.84 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 195.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 190.235 18.96 190.565 ;
      VIA 18.17 190.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 190.215 18.94 190.585 ;
      VIA 18.17 190.4 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 190.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 184.795 18.96 185.125 ;
      VIA 18.17 184.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 184.775 18.94 185.145 ;
      VIA 18.17 184.96 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 184.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 179.355 18.96 179.685 ;
      VIA 18.17 179.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 179.335 18.94 179.705 ;
      VIA 18.17 179.52 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 179.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 173.915 18.96 174.245 ;
      VIA 18.17 174.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 173.895 18.94 174.265 ;
      VIA 18.17 174.08 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 174.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 168.475 18.96 168.805 ;
      VIA 18.17 168.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 168.455 18.94 168.825 ;
      VIA 18.17 168.64 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 168.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 163.035 18.96 163.365 ;
      VIA 18.17 163.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 163.015 18.94 163.385 ;
      VIA 18.17 163.2 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 163.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 157.595 18.96 157.925 ;
      VIA 18.17 157.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 157.575 18.94 157.945 ;
      VIA 18.17 157.76 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 157.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 152.155 18.96 152.485 ;
      VIA 18.17 152.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 152.135 18.94 152.505 ;
      VIA 18.17 152.32 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 152.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 146.715 18.96 147.045 ;
      VIA 18.17 146.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 146.695 18.94 147.065 ;
      VIA 18.17 146.88 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 146.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 141.275 18.96 141.605 ;
      VIA 18.17 141.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 141.255 18.94 141.625 ;
      VIA 18.17 141.44 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 141.44 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 135.835 18.96 136.165 ;
      VIA 18.17 136 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 135.815 18.94 136.185 ;
      VIA 18.17 136 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 136 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 130.395 18.96 130.725 ;
      VIA 18.17 130.56 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 130.375 18.94 130.745 ;
      VIA 18.17 130.56 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 130.56 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 124.955 18.96 125.285 ;
      VIA 18.17 125.12 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 124.935 18.94 125.305 ;
      VIA 18.17 125.12 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 125.12 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 119.515 18.96 119.845 ;
      VIA 18.17 119.68 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 119.495 18.94 119.865 ;
      VIA 18.17 119.68 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 119.68 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 114.075 18.96 114.405 ;
      VIA 18.17 114.24 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 114.055 18.94 114.425 ;
      VIA 18.17 114.24 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 114.24 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 108.635 18.96 108.965 ;
      VIA 18.17 108.8 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 108.615 18.94 108.985 ;
      VIA 18.17 108.8 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 108.8 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 103.195 18.96 103.525 ;
      VIA 18.17 103.36 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 103.175 18.94 103.545 ;
      VIA 18.17 103.36 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 103.36 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 97.755 18.96 98.085 ;
      VIA 18.17 97.92 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 97.735 18.94 98.105 ;
      VIA 18.17 97.92 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 97.92 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 92.315 18.96 92.645 ;
      VIA 18.17 92.48 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 92.295 18.94 92.665 ;
      VIA 18.17 92.48 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 92.48 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 86.875 18.96 87.205 ;
      VIA 18.17 87.04 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 86.855 18.94 87.225 ;
      VIA 18.17 87.04 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 87.04 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 81.435 18.96 81.765 ;
      VIA 18.17 81.6 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 81.415 18.94 81.785 ;
      VIA 18.17 81.6 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 81.6 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 75.995 18.96 76.325 ;
      VIA 18.17 76.16 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 75.975 18.94 76.345 ;
      VIA 18.17 76.16 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 76.16 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 70.555 18.96 70.885 ;
      VIA 18.17 70.72 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 70.535 18.94 70.905 ;
      VIA 18.17 70.72 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 70.72 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 65.115 18.96 65.445 ;
      VIA 18.17 65.28 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 65.095 18.94 65.465 ;
      VIA 18.17 65.28 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 65.28 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 59.675 18.96 60.005 ;
      VIA 18.17 59.84 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 59.655 18.94 60.025 ;
      VIA 18.17 59.84 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 59.84 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 54.235 18.96 54.565 ;
      VIA 18.17 54.4 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 54.215 18.94 54.585 ;
      VIA 18.17 54.4 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 54.4 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 48.795 18.96 49.125 ;
      VIA 18.17 48.96 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 48.775 18.94 49.145 ;
      VIA 18.17 48.96 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 48.96 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 43.355 18.96 43.685 ;
      VIA 18.17 43.52 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 43.335 18.94 43.705 ;
      VIA 18.17 43.52 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 43.52 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 37.915 18.96 38.245 ;
      VIA 18.17 38.08 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 37.895 18.94 38.265 ;
      VIA 18.17 38.08 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 38.08 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 32.475 18.96 32.805 ;
      VIA 18.17 32.64 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 32.455 18.94 32.825 ;
      VIA 18.17 32.64 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 32.64 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 27.035 18.96 27.365 ;
      VIA 18.17 27.2 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 27.015 18.94 27.385 ;
      VIA 18.17 27.2 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 27.2 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 21.595 18.96 21.925 ;
      VIA 18.17 21.76 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 21.575 18.94 21.945 ;
      VIA 18.17 21.76 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 21.76 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 16.155 18.96 16.485 ;
      VIA 18.17 16.32 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 16.135 18.94 16.505 ;
      VIA 18.17 16.32 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 16.32 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 10.715 18.96 11.045 ;
      VIA 18.17 10.88 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 10.695 18.94 11.065 ;
      VIA 18.17 10.88 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 10.88 via2_3_1600_480_1_5_320_320 ;
      LAYER met3 ;
        RECT  17.38 5.275 18.96 5.605 ;
      VIA 18.17 5.44 via4_5_1600_480_1_4_400_400 ;
      LAYER met2 ;
        RECT  17.4 5.255 18.94 5.625 ;
      VIA 18.17 5.44 via3_4_1600_480_1_4_400_400 ;
      VIA 18.17 5.44 via2_3_1600_480_1_5_320_320 ;
    END
  END VSS
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  274.32 288.4 274.46 288.885 ;
    END
  END clk
  PIN i_dbus_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 12.43 288.885 12.73 ;
    END
  END i_dbus_ack
  PIN i_dbus_rdt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  87.56 288.4 87.7 288.885 ;
    END
  END i_dbus_rdt[0]
  PIN i_dbus_rdt[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  84.8 288.4 84.94 288.885 ;
    END
  END i_dbus_rdt[10]
  PIN i_dbus_rdt[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 190.59 0.8 190.89 ;
    END
  END i_dbus_rdt[11]
  PIN i_dbus_rdt[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  105.04 0 105.18 0.485 ;
    END
  END i_dbus_rdt[12]
  PIN i_dbus_rdt[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  233.84 0 233.98 0.485 ;
    END
  END i_dbus_rdt[13]
  PIN i_dbus_rdt[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  276.16 0 276.3 0.485 ;
    END
  END i_dbus_rdt[14]
  PIN i_dbus_rdt[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  277.08 0 277.22 0.485 ;
    END
  END i_dbus_rdt[15]
  PIN i_dbus_rdt[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 99.47 288.885 99.77 ;
    END
  END i_dbus_rdt[16]
  PIN i_dbus_rdt[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 104.91 288.885 105.21 ;
    END
  END i_dbus_rdt[17]
  PIN i_dbus_rdt[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  140.92 0 141.06 0.485 ;
    END
  END i_dbus_rdt[18]
  PIN i_dbus_rdt[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.52 0 99.66 0.485 ;
    END
  END i_dbus_rdt[19]
  PIN i_dbus_rdt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  88.48 0 88.62 0.485 ;
    END
  END i_dbus_rdt[1]
  PIN i_dbus_rdt[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  96.76 288.4 96.9 288.885 ;
    END
  END i_dbus_rdt[20]
  PIN i_dbus_rdt[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  243.96 0 244.1 0.485 ;
    END
  END i_dbus_rdt[21]
  PIN i_dbus_rdt[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  142.76 0 142.9 0.485 ;
    END
  END i_dbus_rdt[22]
  PIN i_dbus_rdt[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  136.32 288.4 136.46 288.885 ;
    END
  END i_dbus_rdt[23]
  PIN i_dbus_rdt[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 98.11 288.885 98.41 ;
    END
  END i_dbus_rdt[24]
  PIN i_dbus_rdt[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 96.75 288.885 97.05 ;
    END
  END i_dbus_rdt[25]
  PIN i_dbus_rdt[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  67.32 0 67.46 0.485 ;
    END
  END i_dbus_rdt[26]
  PIN i_dbus_rdt[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  226.48 0 226.62 0.485 ;
    END
  END i_dbus_rdt[27]
  PIN i_dbus_rdt[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  186.92 0 187.06 0.485 ;
    END
  END i_dbus_rdt[28]
  PIN i_dbus_rdt[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 79.07 288.885 79.37 ;
    END
  END i_dbus_rdt[29]
  PIN i_dbus_rdt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 149.79 0.8 150.09 ;
    END
  END i_dbus_rdt[2]
  PIN i_dbus_rdt[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 178.35 288.885 178.65 ;
    END
  END i_dbus_rdt[30]
  PIN i_dbus_rdt[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  94.92 288.4 95.06 288.885 ;
    END
  END i_dbus_rdt[31]
  PIN i_dbus_rdt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.76 288.4 73.9 288.885 ;
    END
  END i_dbus_rdt[3]
  PIN i_dbus_rdt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 172.91 0.8 173.21 ;
    END
  END i_dbus_rdt[4]
  PIN i_dbus_rdt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 159.31 0.8 159.61 ;
    END
  END i_dbus_rdt[5]
  PIN i_dbus_rdt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  164.84 288.4 164.98 288.885 ;
    END
  END i_dbus_rdt[6]
  PIN i_dbus_rdt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 273.55 288.885 273.85 ;
    END
  END i_dbus_rdt[7]
  PIN i_dbus_rdt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  100.44 0 100.58 0.485 ;
    END
  END i_dbus_rdt[8]
  PIN i_dbus_rdt[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  94 288.4 94.14 288.885 ;
    END
  END i_dbus_rdt[9]
  PIN i_ext_rd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  1.08 0 1.22 0.485 ;
    END
  END i_ext_rd[0]
  PIN i_ext_rd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2 0 2.14 0.485 ;
    END
  END i_ext_rd[10]
  PIN i_ext_rd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2.92 0 3.06 0.485 ;
    END
  END i_ext_rd[11]
  PIN i_ext_rd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  3.84 0 3.98 0.485 ;
    END
  END i_ext_rd[12]
  PIN i_ext_rd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  4.76 0 4.9 0.485 ;
    END
  END i_ext_rd[13]
  PIN i_ext_rd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  5.68 0 5.82 0.485 ;
    END
  END i_ext_rd[14]
  PIN i_ext_rd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  6.6 0 6.74 0.485 ;
    END
  END i_ext_rd[15]
  PIN i_ext_rd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  7.52 0 7.66 0.485 ;
    END
  END i_ext_rd[16]
  PIN i_ext_rd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  8.44 0 8.58 0.485 ;
    END
  END i_ext_rd[17]
  PIN i_ext_rd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  9.36 0 9.5 0.485 ;
    END
  END i_ext_rd[18]
  PIN i_ext_rd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  10.28 0 10.42 0.485 ;
    END
  END i_ext_rd[19]
  PIN i_ext_rd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  11.2 0 11.34 0.485 ;
    END
  END i_ext_rd[1]
  PIN i_ext_rd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  12.12 0 12.26 0.485 ;
    END
  END i_ext_rd[20]
  PIN i_ext_rd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.04 0 13.18 0.485 ;
    END
  END i_ext_rd[21]
  PIN i_ext_rd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  13.96 0 14.1 0.485 ;
    END
  END i_ext_rd[22]
  PIN i_ext_rd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  14.88 0 15.02 0.485 ;
    END
  END i_ext_rd[23]
  PIN i_ext_rd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  15.8 0 15.94 0.485 ;
    END
  END i_ext_rd[24]
  PIN i_ext_rd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  16.72 0 16.86 0.485 ;
    END
  END i_ext_rd[25]
  PIN i_ext_rd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  17.64 0 17.78 0.485 ;
    END
  END i_ext_rd[26]
  PIN i_ext_rd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  18.56 0 18.7 0.485 ;
    END
  END i_ext_rd[27]
  PIN i_ext_rd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  19.48 0 19.62 0.485 ;
    END
  END i_ext_rd[28]
  PIN i_ext_rd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  20.4 0 20.54 0.485 ;
    END
  END i_ext_rd[29]
  PIN i_ext_rd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  21.32 0 21.46 0.485 ;
    END
  END i_ext_rd[2]
  PIN i_ext_rd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  22.24 0 22.38 0.485 ;
    END
  END i_ext_rd[30]
  PIN i_ext_rd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  23.16 0 23.3 0.485 ;
    END
  END i_ext_rd[31]
  PIN i_ext_rd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  24.08 0 24.22 0.485 ;
    END
  END i_ext_rd[3]
  PIN i_ext_rd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25 0 25.14 0.485 ;
    END
  END i_ext_rd[4]
  PIN i_ext_rd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  25.92 0 26.06 0.485 ;
    END
  END i_ext_rd[5]
  PIN i_ext_rd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  26.84 0 26.98 0.485 ;
    END
  END i_ext_rd[6]
  PIN i_ext_rd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  27.76 0 27.9 0.485 ;
    END
  END i_ext_rd[7]
  PIN i_ext_rd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  28.68 0 28.82 0.485 ;
    END
  END i_ext_rd[8]
  PIN i_ext_rd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  29.6 0 29.74 0.485 ;
    END
  END i_ext_rd[9]
  PIN i_ext_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  30.52 0 30.66 0.485 ;
    END
  END i_ext_ready
  PIN i_ibus_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 259.95 0.8 260.25 ;
    END
  END i_ibus_ack
  PIN i_ibus_rdt[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  31.44 0 31.58 0.485 ;
    END
  END i_ibus_rdt[0]
  PIN i_ibus_rdt[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  197.96 288.4 198.1 288.885 ;
    END
  END i_ibus_rdt[10]
  PIN i_ibus_rdt[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  196.12 288.4 196.26 288.885 ;
    END
  END i_ibus_rdt[11]
  PIN i_ibus_rdt[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 142.99 0.8 143.29 ;
    END
  END i_ibus_rdt[12]
  PIN i_ibus_rdt[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 142.99 288.885 143.29 ;
    END
  END i_ibus_rdt[13]
  PIN i_ibus_rdt[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 164.75 0.8 165.05 ;
    END
  END i_ibus_rdt[14]
  PIN i_ibus_rdt[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  143.68 0 143.82 0.485 ;
    END
  END i_ibus_rdt[15]
  PIN i_ibus_rdt[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 111.71 288.885 112.01 ;
    END
  END i_ibus_rdt[16]
  PIN i_ibus_rdt[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  153.8 288.4 153.94 288.885 ;
    END
  END i_ibus_rdt[17]
  PIN i_ibus_rdt[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  145.52 288.4 145.66 288.885 ;
    END
  END i_ibus_rdt[18]
  PIN i_ibus_rdt[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  138.16 288.4 138.3 288.885 ;
    END
  END i_ibus_rdt[19]
  PIN i_ibus_rdt[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  32.36 0 32.5 0.485 ;
    END
  END i_ibus_rdt[1]
  PIN i_ibus_rdt[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  150.12 288.4 150.26 288.885 ;
    END
  END i_ibus_rdt[20]
  PIN i_ibus_rdt[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  147.36 288.4 147.5 288.885 ;
    END
  END i_ibus_rdt[21]
  PIN i_ibus_rdt[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  163 288.4 163.14 288.885 ;
    END
  END i_ibus_rdt[22]
  PIN i_ibus_rdt[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  101.36 288.4 101.5 288.885 ;
    END
  END i_ibus_rdt[23]
  PIN i_ibus_rdt[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  99.52 288.4 99.66 288.885 ;
    END
  END i_ibus_rdt[24]
  PIN i_ibus_rdt[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  174.96 288.4 175.1 288.885 ;
    END
  END i_ibus_rdt[25]
  PIN i_ibus_rdt[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  163.92 288.4 164.06 288.885 ;
    END
  END i_ibus_rdt[26]
  PIN i_ibus_rdt[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  102.28 288.4 102.42 288.885 ;
    END
  END i_ibus_rdt[27]
  PIN i_ibus_rdt[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 152.51 0.8 152.81 ;
    END
  END i_ibus_rdt[28]
  PIN i_ibus_rdt[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 137.55 0.8 137.85 ;
    END
  END i_ibus_rdt[29]
  PIN i_ibus_rdt[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 182.43 0.8 182.73 ;
    END
  END i_ibus_rdt[2]
  PIN i_ibus_rdt[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 136.19 0.8 136.49 ;
    END
  END i_ibus_rdt[30]
  PIN i_ibus_rdt[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  90.32 288.4 90.46 288.885 ;
    END
  END i_ibus_rdt[31]
  PIN i_ibus_rdt[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  98.6 288.4 98.74 288.885 ;
    END
  END i_ibus_rdt[3]
  PIN i_ibus_rdt[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  97.68 288.4 97.82 288.885 ;
    END
  END i_ibus_rdt[4]
  PIN i_ibus_rdt[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 230.03 0.8 230.33 ;
    END
  END i_ibus_rdt[5]
  PIN i_ibus_rdt[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 186.51 0.8 186.81 ;
    END
  END i_ibus_rdt[6]
  PIN i_ibus_rdt[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  199.8 288.4 199.94 288.885 ;
    END
  END i_ibus_rdt[7]
  PIN i_ibus_rdt[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  206.24 288.4 206.38 288.885 ;
    END
  END i_ibus_rdt[8]
  PIN i_ibus_rdt[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  204.4 288.4 204.54 288.885 ;
    END
  END i_ibus_rdt[9]
  PIN i_rdata0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 212.35 0.8 212.65 ;
    END
  END i_rdata0
  PIN i_rdata1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  169.44 288.4 169.58 288.885 ;
    END
  END i_rdata1
  PIN i_rf_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  191.52 288.4 191.66 288.885 ;
    END
  END i_rf_ready
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  202.56 288.4 202.7 288.885 ;
    END
  END i_rst
  PIN i_timer_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  187.84 288.4 187.98 288.885 ;
    END
  END i_timer_irq
  PIN o_dbus_adr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 276.27 0.8 276.57 ;
    END
  END o_dbus_adr[0]
  PIN o_dbus_adr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  196.12 0 196.26 0.485 ;
    END
  END o_dbus_adr[10]
  PIN o_dbus_adr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 68.19 288.885 68.49 ;
    END
  END o_dbus_adr[11]
  PIN o_dbus_adr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 274.91 288.885 275.21 ;
    END
  END o_dbus_adr[12]
  PIN o_dbus_adr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 36.91 288.885 37.21 ;
    END
  END o_dbus_adr[13]
  PIN o_dbus_adr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  209.92 0 210.06 0.485 ;
    END
  END o_dbus_adr[14]
  PIN o_dbus_adr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 114.43 288.885 114.73 ;
    END
  END o_dbus_adr[15]
  PIN o_dbus_adr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  225.56 0 225.7 0.485 ;
    END
  END o_dbus_adr[16]
  PIN o_dbus_adr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 128.03 0.8 128.33 ;
    END
  END o_dbus_adr[17]
  PIN o_dbus_adr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  188.76 0 188.9 0.485 ;
    END
  END o_dbus_adr[18]
  PIN o_dbus_adr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  190.6 0 190.74 0.485 ;
    END
  END o_dbus_adr[19]
  PIN o_dbus_adr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 5.63 0.8 5.93 ;
    END
  END o_dbus_adr[1]
  PIN o_dbus_adr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 65.47 288.885 65.77 ;
    END
  END o_dbus_adr[20]
  PIN o_dbus_adr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  189.68 0 189.82 0.485 ;
    END
  END o_dbus_adr[21]
  PIN o_dbus_adr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  109.64 0 109.78 0.485 ;
    END
  END o_dbus_adr[22]
  PIN o_dbus_adr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  193.36 0 193.5 0.485 ;
    END
  END o_dbus_adr[23]
  PIN o_dbus_adr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  206.24 0 206.38 0.485 ;
    END
  END o_dbus_adr[24]
  PIN o_dbus_adr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  207.16 0 207.3 0.485 ;
    END
  END o_dbus_adr[25]
  PIN o_dbus_adr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  271.56 288.4 271.7 288.885 ;
    END
  END o_dbus_adr[26]
  PIN o_dbus_adr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  186 288.4 186.14 288.885 ;
    END
  END o_dbus_adr[27]
  PIN o_dbus_adr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  183.24 288.4 183.38 288.885 ;
    END
  END o_dbus_adr[28]
  PIN o_dbus_adr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 270.83 0.8 271.13 ;
    END
  END o_dbus_adr[29]
  PIN o_dbus_adr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 145.71 288.885 146.01 ;
    END
  END o_dbus_adr[2]
  PIN o_dbus_adr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  89.4 288.4 89.54 288.885 ;
    END
  END o_dbus_adr[30]
  PIN o_dbus_adr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 113.07 288.885 113.37 ;
    END
  END o_dbus_adr[31]
  PIN o_dbus_adr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 281.71 288.885 282.01 ;
    END
  END o_dbus_adr[3]
  PIN o_dbus_adr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 280.35 288.885 280.65 ;
    END
  END o_dbus_adr[4]
  PIN o_dbus_adr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  222.8 288.4 222.94 288.885 ;
    END
  END o_dbus_adr[5]
  PIN o_dbus_adr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  80.2 288.4 80.34 288.885 ;
    END
  END o_dbus_adr[6]
  PIN o_dbus_adr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  85.72 288.4 85.86 288.885 ;
    END
  END o_dbus_adr[7]
  PIN o_dbus_adr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 122.59 288.885 122.89 ;
    END
  END o_dbus_adr[8]
  PIN o_dbus_adr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  123.44 0 123.58 0.485 ;
    END
  END o_dbus_adr[9]
  PIN o_dbus_cyc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 167.47 0.8 167.77 ;
    END
  END o_dbus_cyc
  PIN o_dbus_dat[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  81.12 0 81.26 0.485 ;
    END
  END o_dbus_dat[0]
  PIN o_dbus_dat[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  88.48 288.4 88.62 288.885 ;
    END
  END o_dbus_dat[10]
  PIN o_dbus_dat[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 273.55 0.8 273.85 ;
    END
  END o_dbus_dat[11]
  PIN o_dbus_dat[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  66.4 0 66.54 0.485 ;
    END
  END o_dbus_dat[12]
  PIN o_dbus_dat[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  33.28 0 33.42 0.485 ;
    END
  END o_dbus_dat[13]
  PIN o_dbus_dat[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  234.76 0 234.9 0.485 ;
    END
  END o_dbus_dat[14]
  PIN o_dbus_dat[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  209 0 209.14 0.485 ;
    END
  END o_dbus_dat[15]
  PIN o_dbus_dat[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 13.79 288.885 14.09 ;
    END
  END o_dbus_dat[16]
  PIN o_dbus_dat[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  187.84 0 187.98 0.485 ;
    END
  END o_dbus_dat[17]
  PIN o_dbus_dat[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  165.76 288.4 165.9 288.885 ;
    END
  END o_dbus_dat[18]
  PIN o_dbus_dat[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  101.36 0 101.5 0.485 ;
    END
  END o_dbus_dat[19]
  PIN o_dbus_dat[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  34.2 0 34.34 0.485 ;
    END
  END o_dbus_dat[1]
  PIN o_dbus_dat[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  184.16 288.4 184.3 288.885 ;
    END
  END o_dbus_dat[20]
  PIN o_dbus_dat[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 19.23 288.885 19.53 ;
    END
  END o_dbus_dat[21]
  PIN o_dbus_dat[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  199.8 0 199.94 0.485 ;
    END
  END o_dbus_dat[22]
  PIN o_dbus_dat[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  134.48 0 134.62 0.485 ;
    END
  END o_dbus_dat[23]
  PIN o_dbus_dat[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 117.15 288.885 117.45 ;
    END
  END o_dbus_dat[24]
  PIN o_dbus_dat[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 95.39 288.885 95.69 ;
    END
  END o_dbus_dat[25]
  PIN o_dbus_dat[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  35.12 0 35.26 0.485 ;
    END
  END o_dbus_dat[26]
  PIN o_dbus_dat[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  36.04 0 36.18 0.485 ;
    END
  END o_dbus_dat[27]
  PIN o_dbus_dat[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  203.48 0 203.62 0.485 ;
    END
  END o_dbus_dat[28]
  PIN o_dbus_dat[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  73.76 0 73.9 0.485 ;
    END
  END o_dbus_dat[29]
  PIN o_dbus_dat[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  86.64 288.4 86.78 288.885 ;
    END
  END o_dbus_dat[2]
  PIN o_dbus_dat[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  223.72 0 223.86 0.485 ;
    END
  END o_dbus_dat[30]
  PIN o_dbus_dat[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  201.64 0 201.78 0.485 ;
    END
  END o_dbus_dat[31]
  PIN o_dbus_dat[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  91.24 288.4 91.38 288.885 ;
    END
  END o_dbus_dat[3]
  PIN o_dbus_dat[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 171.55 288.885 171.85 ;
    END
  END o_dbus_dat[4]
  PIN o_dbus_dat[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 176.99 0.8 177.29 ;
    END
  END o_dbus_dat[5]
  PIN o_dbus_dat[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  93.08 288.4 93.22 288.885 ;
    END
  END o_dbus_dat[6]
  PIN o_dbus_dat[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  248.56 288.4 248.7 288.885 ;
    END
  END o_dbus_dat[7]
  PIN o_dbus_dat[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 208.27 0.8 208.57 ;
    END
  END o_dbus_dat[8]
  PIN o_dbus_dat[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  47.08 0 47.22 0.485 ;
    END
  END o_dbus_dat[9]
  PIN o_dbus_sel[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  89.4 0 89.54 0.485 ;
    END
  END o_dbus_sel[0]
  PIN o_dbus_sel[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 147.07 0.8 147.37 ;
    END
  END o_dbus_sel[1]
  PIN o_dbus_sel[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  108.72 0 108.86 0.485 ;
    END
  END o_dbus_sel[2]
  PIN o_dbus_sel[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 141.63 0.8 141.93 ;
    END
  END o_dbus_sel[3]
  PIN o_dbus_we
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  149.2 288.4 149.34 288.885 ;
    END
  END o_dbus_we
  PIN o_ext_funct3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 200.11 0.8 200.41 ;
    END
  END o_ext_funct3[0]
  PIN o_ext_funct3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 80.43 288.885 80.73 ;
    END
  END o_ext_funct3[1]
  PIN o_ext_funct3[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 224.59 0.8 224.89 ;
    END
  END o_ext_funct3[2]
  PIN o_ext_rs1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  90.32 0 90.46 0.485 ;
    END
  END o_ext_rs1[0]
  PIN o_ext_rs1[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  202.56 0 202.7 0.485 ;
    END
  END o_ext_rs1[10]
  PIN o_ext_rs1[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 69.55 288.885 69.85 ;
    END
  END o_ext_rs1[11]
  PIN o_ext_rs1[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 276.27 288.885 276.57 ;
    END
  END o_ext_rs1[12]
  PIN o_ext_rs1[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  278.92 0 279.06 0.485 ;
    END
  END o_ext_rs1[13]
  PIN o_ext_rs1[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  155.64 0 155.78 0.485 ;
    END
  END o_ext_rs1[14]
  PIN o_ext_rs1[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 272.19 288.885 272.49 ;
    END
  END o_ext_rs1[15]
  PIN o_ext_rs1[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  228.32 0 228.46 0.485 ;
    END
  END o_ext_rs1[16]
  PIN o_ext_rs1[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 129.39 0.8 129.69 ;
    END
  END o_ext_rs1[17]
  PIN o_ext_rs1[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  191.52 0 191.66 0.485 ;
    END
  END o_ext_rs1[18]
  PIN o_ext_rs1[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  195.2 0 195.34 0.485 ;
    END
  END o_ext_rs1[19]
  PIN o_ext_rs1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  91.24 0 91.38 0.485 ;
    END
  END o_ext_rs1[1]
  PIN o_ext_rs1[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 64.11 288.885 64.41 ;
    END
  END o_ext_rs1[20]
  PIN o_ext_rs1[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  121.6 0 121.74 0.485 ;
    END
  END o_ext_rs1[21]
  PIN o_ext_rs1[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  107.8 0 107.94 0.485 ;
    END
  END o_ext_rs1[22]
  PIN o_ext_rs1[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  194.28 0 194.42 0.485 ;
    END
  END o_ext_rs1[23]
  PIN o_ext_rs1[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  205.32 0 205.46 0.485 ;
    END
  END o_ext_rs1[24]
  PIN o_ext_rs1[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  208.08 0 208.22 0.485 ;
    END
  END o_ext_rs1[25]
  PIN o_ext_rs1[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  95.84 288.4 95.98 288.885 ;
    END
  END o_ext_rs1[26]
  PIN o_ext_rs1[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  103.2 288.4 103.34 288.885 ;
    END
  END o_ext_rs1[27]
  PIN o_ext_rs1[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  185.08 288.4 185.22 288.885 ;
    END
  END o_ext_rs1[28]
  PIN o_ext_rs1[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 13.79 0.8 14.09 ;
    END
  END o_ext_rs1[29]
  PIN o_ext_rs1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 144.35 288.885 144.65 ;
    END
  END o_ext_rs1[2]
  PIN o_ext_rs1[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  170.36 288.4 170.5 288.885 ;
    END
  END o_ext_rs1[30]
  PIN o_ext_rs1[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 106.27 288.885 106.57 ;
    END
  END o_ext_rs1[31]
  PIN o_ext_rs1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 278.99 288.885 279.29 ;
    END
  END o_ext_rs1[3]
  PIN o_ext_rs1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  227.4 288.4 227.54 288.885 ;
    END
  END o_ext_rs1[4]
  PIN o_ext_rs1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  142.76 288.4 142.9 288.885 ;
    END
  END o_ext_rs1[5]
  PIN o_ext_rs1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  10.28 288.4 10.42 288.885 ;
    END
  END o_ext_rs1[6]
  PIN o_ext_rs1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  78.36 288.4 78.5 288.885 ;
    END
  END o_ext_rs1[7]
  PIN o_ext_rs1[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 123.95 288.885 124.25 ;
    END
  END o_ext_rs1[8]
  PIN o_ext_rs1[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  122.52 0 122.66 0.485 ;
    END
  END o_ext_rs1[9]
  PIN o_ext_rs2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  136.32 0 136.46 0.485 ;
    END
  END o_ext_rs2[0]
  PIN o_ext_rs2[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  66.4 288.4 66.54 288.885 ;
    END
  END o_ext_rs2[10]
  PIN o_ext_rs2[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 115.79 0.8 116.09 ;
    END
  END o_ext_rs2[11]
  PIN o_ext_rs2[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  204.4 0 204.54 0.485 ;
    END
  END o_ext_rs2[12]
  PIN o_ext_rs2[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 16.51 0.8 16.81 ;
    END
  END o_ext_rs2[13]
  PIN o_ext_rs2[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 51.87 288.885 52.17 ;
    END
  END o_ext_rs2[14]
  PIN o_ext_rs2[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  128.04 0 128.18 0.485 ;
    END
  END o_ext_rs2[15]
  PIN o_ext_rs2[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  185.08 0 185.22 0.485 ;
    END
  END o_ext_rs2[16]
  PIN o_ext_rs2[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  268.8 0 268.94 0.485 ;
    END
  END o_ext_rs2[17]
  PIN o_ext_rs2[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  141.84 288.4 141.98 288.885 ;
    END
  END o_ext_rs2[18]
  PIN o_ext_rs2[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  120.68 0 120.82 0.485 ;
    END
  END o_ext_rs2[19]
  PIN o_ext_rs2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 6.99 0.8 7.29 ;
    END
  END o_ext_rs2[1]
  PIN o_ext_rs2[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  186.92 288.4 187.06 288.885 ;
    END
  END o_ext_rs2[20]
  PIN o_ext_rs2[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 88.59 288.885 88.89 ;
    END
  END o_ext_rs2[21]
  PIN o_ext_rs2[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 94.03 288.885 94.33 ;
    END
  END o_ext_rs2[22]
  PIN o_ext_rs2[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  135.4 0 135.54 0.485 ;
    END
  END o_ext_rs2[23]
  PIN o_ext_rs2[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 277.63 288.885 277.93 ;
    END
  END o_ext_rs2[24]
  PIN o_ext_rs2[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 92.67 288.885 92.97 ;
    END
  END o_ext_rs2[25]
  PIN o_ext_rs2[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 15.15 0.8 15.45 ;
    END
  END o_ext_rs2[26]
  PIN o_ext_rs2[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 96.75 0.8 97.05 ;
    END
  END o_ext_rs2[27]
  PIN o_ext_rs2[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  186 0 186.14 0.485 ;
    END
  END o_ext_rs2[28]
  PIN o_ext_rs2[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  74.68 0 74.82 0.485 ;
    END
  END o_ext_rs2[29]
  PIN o_ext_rs2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  77.44 288.4 77.58 288.885 ;
    END
  END o_ext_rs2[2]
  PIN o_ext_rs2[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  224.64 0 224.78 0.485 ;
    END
  END o_ext_rs2[30]
  PIN o_ext_rs2[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  278 0 278.14 0.485 ;
    END
  END o_ext_rs2[31]
  PIN o_ext_rs2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  100.44 288.4 100.58 288.885 ;
    END
  END o_ext_rs2[3]
  PIN o_ext_rs2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 194.67 288.885 194.97 ;
    END
  END o_ext_rs2[4]
  PIN o_ext_rs2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 178.35 0.8 178.65 ;
    END
  END o_ext_rs2[5]
  PIN o_ext_rs2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  64.56 288.4 64.7 288.885 ;
    END
  END o_ext_rs2[6]
  PIN o_ext_rs2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  158.4 288.4 158.54 288.885 ;
    END
  END o_ext_rs2[7]
  PIN o_ext_rs2[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 11.07 0.8 11.37 ;
    END
  END o_ext_rs2[8]
  PIN o_ext_rs2[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 8.35 0.8 8.65 ;
    END
  END o_ext_rs2[9]
  PIN o_ibus_adr[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 91.31 288.885 91.61 ;
    END
  END o_ibus_adr[0]
  PIN o_ibus_adr[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 89.95 288.885 90.25 ;
    END
  END o_ibus_adr[10]
  PIN o_ibus_adr[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 152.51 288.885 152.81 ;
    END
  END o_ibus_adr[11]
  PIN o_ibus_adr[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 159.31 288.885 159.61 ;
    END
  END o_ibus_adr[12]
  PIN o_ibus_adr[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 166.11 288.885 166.41 ;
    END
  END o_ibus_adr[13]
  PIN o_ibus_adr[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 164.75 288.885 165.05 ;
    END
  END o_ibus_adr[14]
  PIN o_ibus_adr[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 167.47 288.885 167.77 ;
    END
  END o_ibus_adr[15]
  PIN o_ibus_adr[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 175.63 288.885 175.93 ;
    END
  END o_ibus_adr[16]
  PIN o_ibus_adr[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 183.79 288.885 184.09 ;
    END
  END o_ibus_adr[17]
  PIN o_ibus_adr[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 181.07 288.885 181.37 ;
    END
  END o_ibus_adr[18]
  PIN o_ibus_adr[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 179.71 288.885 180.01 ;
    END
  END o_ibus_adr[19]
  PIN o_ibus_adr[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  235.68 0 235.82 0.485 ;
    END
  END o_ibus_adr[1]
  PIN o_ibus_adr[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 182.43 288.885 182.73 ;
    END
  END o_ibus_adr[20]
  PIN o_ibus_adr[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 121.23 288.885 121.53 ;
    END
  END o_ibus_adr[21]
  PIN o_ibus_adr[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 118.51 288.885 118.81 ;
    END
  END o_ibus_adr[22]
  PIN o_ibus_adr[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 84.51 288.885 84.81 ;
    END
  END o_ibus_adr[23]
  PIN o_ibus_adr[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  198.88 0 199.02 0.485 ;
    END
  END o_ibus_adr[24]
  PIN o_ibus_adr[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  197.04 0 197.18 0.485 ;
    END
  END o_ibus_adr[25]
  PIN o_ibus_adr[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  197.96 0 198.1 0.485 ;
    END
  END o_ibus_adr[26]
  PIN o_ibus_adr[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  200.72 0 200.86 0.485 ;
    END
  END o_ibus_adr[27]
  PIN o_ibus_adr[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  192.44 0 192.58 0.485 ;
    END
  END o_ibus_adr[28]
  PIN o_ibus_adr[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 66.83 288.885 67.13 ;
    END
  END o_ibus_adr[29]
  PIN o_ibus_adr[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  236.6 0 236.74 0.485 ;
    END
  END o_ibus_adr[2]
  PIN o_ibus_adr[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 176.99 288.885 177.29 ;
    END
  END o_ibus_adr[30]
  PIN o_ibus_adr[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 186.51 288.885 186.81 ;
    END
  END o_ibus_adr[31]
  PIN o_ibus_adr[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  241.2 0 241.34 0.485 ;
    END
  END o_ibus_adr[3]
  PIN o_ibus_adr[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  238.44 0 238.58 0.485 ;
    END
  END o_ibus_adr[4]
  PIN o_ibus_adr[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 108.99 288.885 109.29 ;
    END
  END o_ibus_adr[5]
  PIN o_ibus_adr[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 115.79 288.885 116.09 ;
    END
  END o_ibus_adr[6]
  PIN o_ibus_adr[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 162.03 288.885 162.33 ;
    END
  END o_ibus_adr[7]
  PIN o_ibus_adr[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 100.83 288.885 101.13 ;
    END
  END o_ibus_adr[8]
  PIN o_ibus_adr[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  229.24 0 229.38 0.485 ;
    END
  END o_ibus_adr[9]
  PIN o_ibus_cyc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  203.48 288.4 203.62 288.885 ;
    END
  END o_ibus_cyc
  PIN o_mdu_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 134.83 0.8 135.13 ;
    END
  END o_mdu_valid
  PIN o_rf_rreq
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 163.39 0.8 163.69 ;
    END
  END o_rf_rreq
  PIN o_rf_wreq
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 166.11 0.8 166.41 ;
    END
  END o_rf_wreq
  PIN o_rreg0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 162.03 0.8 162.33 ;
    END
  END o_rreg0[0]
  PIN o_rreg0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 110.35 288.885 110.65 ;
    END
  END o_rreg0[1]
  PIN o_rreg0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  155.64 288.4 155.78 288.885 ;
    END
  END o_rreg0[2]
  PIN o_rreg0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  151.04 288.4 151.18 288.885 ;
    END
  END o_rreg0[3]
  PIN o_rreg0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  140 288.4 140.14 288.885 ;
    END
  END o_rreg0[4]
  PIN o_rreg0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 144.35 0.8 144.65 ;
    END
  END o_rreg0[5]
  PIN o_rreg1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  152.88 288.4 153.02 288.885 ;
    END
  END o_rreg1[0]
  PIN o_rreg1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  144.6 288.4 144.74 288.885 ;
    END
  END o_rreg1[1]
  PIN o_rreg1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  148.28 288.4 148.42 288.885 ;
    END
  END o_rreg1[2]
  PIN o_rreg1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  131.72 288.4 131.86 288.885 ;
    END
  END o_rreg1[3]
  PIN o_rreg1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  129.88 288.4 130.02 288.885 ;
    END
  END o_rreg1[4]
  PIN o_rreg1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  216.36 288.4 216.5 288.885 ;
    END
  END o_rreg1[5]
  PIN o_wdata0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  143.68 288.4 143.82 288.885 ;
    END
  END o_wdata0
  PIN o_wdata1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  159.32 288.4 159.46 288.885 ;
    END
  END o_wdata1
  PIN o_wen0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  192.44 288.4 192.58 288.885 ;
    END
  END o_wen0
  PIN o_wen1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  92.16 288.4 92.3 288.885 ;
    END
  END o_wen1
  PIN o_wreg0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  139.08 288.4 139.22 288.885 ;
    END
  END o_wreg0[0]
  PIN o_wreg0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  197.04 288.4 197.18 288.885 ;
    END
  END o_wreg0[1]
  PIN o_wreg0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  209 288.4 209.14 288.885 ;
    END
  END o_wreg0[2]
  PIN o_wreg0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  195.2 288.4 195.34 288.885 ;
    END
  END o_wreg0[3]
  PIN o_wreg0[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  205.32 288.4 205.46 288.885 ;
    END
  END o_wreg0[4]
  PIN o_wreg0[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  201.64 288.4 201.78 288.885 ;
    END
  END o_wreg0[5]
  PIN o_wreg1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  151.96 288.4 152.1 288.885 ;
    END
  END o_wreg1[0]
  PIN o_wreg1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  140.92 288.4 141.06 288.885 ;
    END
  END o_wreg1[1]
  PIN o_wreg1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 9.71 0.8 10.01 ;
    END
  END o_wreg1[2]
  PIN o_wreg1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 12.43 0.8 12.73 ;
    END
  END o_wreg1[3]
  PIN o_wreg1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  11.2 288.4 11.34 288.885 ;
    END
  END o_wreg1[4]
  PIN o_wreg1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  288.085 107.63 288.885 107.93 ;
    END
  END o_wreg1[5]
  OBS
    LAYER li1 ;
     RECT  4.6 5.355 284.28 282.965 ;
    LAYER met1 ;
     RECT  4.3 9.28 4.6 9.42 ;
     RECT  4.3 132.7 4.6 142.02 ;
     RECT  3.84 229.6 4.6 229.74 ;
     RECT  4.6 5.2 90.78 283.12 ;
     RECT  90.78 0.44 91.7 283.12 ;
     RECT  91.7 0.44 110.7 288.22 ;
     RECT  110.7 4.86 138.3 288.22 ;
     RECT  138.3 5.2 160.38 288.22 ;
     RECT  160.38 5.2 187.84 283.12 ;
     RECT  187.84 0.44 269.4 283.12 ;
     RECT  269.4 5.2 284.28 283.12 ;
     RECT  284.28 117.74 284.58 117.88 ;
     RECT  284.28 12 287.34 12.48 ;
     RECT  284.28 101.08 287.8 101.22 ;
     RECT  287.34 12.34 288.26 12.48 ;
     RECT  284.28 77.28 288.26 77.42 ;
     RECT  284.28 273.12 288.72 273.26 ;
    LAYER met2 ;
     RECT  101.82 0.27 103.34 0.34 ;
     RECT  66.4 0.34 109.78 0.44 ;
     RECT  185.08 0.34 210.06 1.63 ;
     RECT  66.4 0.44 110.7 4.86 ;
     RECT  120.68 0.34 143.82 4.86 ;
     RECT  33.28 0.34 36.18 5.255 ;
     RECT  47.08 0.34 47.22 5.255 ;
     RECT  155.64 0.34 155.78 5.255 ;
     RECT  185.08 1.63 210.98 5.255 ;
     RECT  268.8 0.34 279.06 5.255 ;
     RECT  17.4 5.255 18.94 6.22 ;
     RECT  7.52 5.71 7.66 6.56 ;
     RECT  180.24 5.255 210.98 6.56 ;
     RECT  261.66 5.255 279.06 6.56 ;
     RECT  17.4 6.22 20.54 7.21 ;
     RECT  7.06 6.56 7.66 7.58 ;
     RECT  17.4 7.21 18.94 7.58 ;
     RECT  33.28 5.255 47.22 7.975 ;
     RECT  66.4 4.86 143.82 7.975 ;
     RECT  172.66 6.56 210.98 7.975 ;
     RECT  223.72 0.34 244.1 7.975 ;
     RECT  7.06 7.58 18.94 8.94 ;
     RECT  6.6 8.94 18.94 9.28 ;
     RECT  166.67 7.975 210.98 9.62 ;
     RECT  220.95 7.975 249.63 9.62 ;
     RECT  4.3 9.28 18.94 11.29 ;
     RECT  261.66 6.56 279.52 12 ;
     RECT  261.66 12 287.34 12.34 ;
     RECT  30.97 7.975 47.22 13.02 ;
     RECT  153.1 5.255 155.78 13.16 ;
     RECT  29.14 13.02 47.22 15.54 ;
     RECT  30.97 15.54 47.22 16.9 ;
     RECT  166.67 9.62 249.63 17.78 ;
     RECT  6.14 11.29 18.94 19.62 ;
     RECT  58.11 7.975 143.82 20.5 ;
     RECT  153.1 13.16 154.64 20.5 ;
     RECT  58.11 20.5 154.64 24.04 ;
     RECT  30.97 16.9 46.08 26.08 ;
     RECT  14.88 19.62 18.94 26.28 ;
     RECT  30.97 26.08 32.51 26.28 ;
     RECT  58.11 24.04 143.82 48.04 ;
     RECT  153.1 24.04 154.64 48.04 ;
     RECT  58.11 48.04 154.64 58.38 ;
     RECT  124.82 58.38 154.64 59.4 ;
     RECT  125.28 59.4 154.64 63.82 ;
     RECT  166.67 17.78 251.92 70.28 ;
     RECT  220.95 70.28 251.92 71.84 ;
     RECT  261.66 12.34 288.26 71.84 ;
     RECT  220.95 71.84 288.26 77.42 ;
     RECT  166.67 70.28 208.92 82.72 ;
     RECT  166.67 82.72 210.52 94.62 ;
     RECT  220.95 77.42 287.8 94.62 ;
     RECT  14.88 26.28 32.51 96.66 ;
     RECT  166.67 94.62 287.8 96.66 ;
     RECT  13.96 96.66 32.51 96.8 ;
     RECT  13.96 96.8 18.94 96.97 ;
     RECT  165.3 96.66 287.8 101.22 ;
     RECT  165.3 101.22 282.74 101.9 ;
     RECT  125.96 63.82 154.64 107.2 ;
     RECT  165.3 101.9 251.46 107.2 ;
     RECT  261.66 101.9 282.74 107.85 ;
     RECT  14.88 96.97 18.94 115.87 ;
     RECT  261.66 107.85 282.28 117.23 ;
     RECT  261.66 117.23 284.58 117.91 ;
     RECT  58.11 58.38 113.93 123.52 ;
     RECT  125.96 107.2 251.46 123.52 ;
     RECT  58.11 123.52 251.46 123.66 ;
     RECT  206.24 123.66 251.46 126.21 ;
     RECT  7.06 115.87 18.94 126.24 ;
     RECT  6.6 126.24 18.94 126.58 ;
     RECT  5.68 126.58 18.94 129.61 ;
     RECT  206.7 126.21 251.46 132.7 ;
     RECT  261.66 117.91 288.72 132.7 ;
     RECT  206.7 132.7 288.72 134.88 ;
     RECT  206.7 134.88 251.46 135.05 ;
     RECT  6.6 129.61 18.94 142.9 ;
     RECT  6.14 142.9 18.94 144.57 ;
     RECT  261.66 134.88 288.72 145.62 ;
     RECT  58.11 123.66 196.72 146.44 ;
     RECT  206.7 135.05 250.54 147.66 ;
     RECT  206.24 147.66 250.54 147.8 ;
     RECT  206.7 147.8 250.54 149.02 ;
     RECT  260.98 145.62 288.72 149.02 ;
     RECT  58.11 146.44 195.35 158.88 ;
     RECT  206.7 149.02 288.72 158.88 ;
     RECT  30.97 96.8 32.51 181.66 ;
     RECT  44.54 26.08 46.08 181.66 ;
     RECT  58.11 158.88 288.72 183.84 ;
     RECT  58.11 183.84 238.12 184.52 ;
     RECT  58.11 184.52 237.66 185.88 ;
     RECT  218.2 185.88 222.94 186.22 ;
     RECT  220.95 186.22 222.94 188.26 ;
     RECT  232.46 185.88 237.66 188.26 ;
     RECT  232.46 188.26 236.06 189.96 ;
     RECT  58.11 185.88 208.92 191.66 ;
     RECT  69.62 191.66 208.92 205.46 ;
     RECT  69.16 205.46 208.92 207.64 ;
     RECT  248.09 183.84 288.72 211.04 ;
     RECT  234.52 189.96 236.06 211.58 ;
     RECT  248.09 211.04 250.54 211.58 ;
     RECT  14.88 144.57 18.94 220.76 ;
     RECT  69.62 207.64 208.92 222.12 ;
     RECT  14.42 220.76 18.94 227.56 ;
     RECT  69.62 222.12 209.6 227.63 ;
     RECT  9.82 227.56 18.94 229.06 ;
     RECT  3.84 229.6 3.98 230.25 ;
     RECT  30.97 181.66 46.08 232.8 ;
     RECT  69.16 227.63 209.6 241.16 ;
     RECT  220.95 188.26 222.49 241.16 ;
     RECT  69.16 241.16 222.49 252.01 ;
     RECT  69.16 252.01 100.36 262.24 ;
     RECT  69.16 262.24 101.96 262.75 ;
     RECT  111.48 252.01 222.49 262.75 ;
     RECT  13.96 229.06 18.94 268.7 ;
     RECT  44.54 232.8 46.08 268.7 ;
     RECT  69.16 262.75 222.49 269.72 ;
     RECT  234.52 211.58 250.54 269.72 ;
     RECT  69.16 269.72 250.54 269.86 ;
     RECT  71.68 269.86 250.54 270.06 ;
     RECT  261.66 211.04 288.72 270.06 ;
     RECT  71.68 270.06 288.72 273.26 ;
     RECT  71.68 273.26 282.74 275.64 ;
     RECT  71.68 275.64 250.08 275.98 ;
     RECT  10.28 268.7 18.94 276.35 ;
     RECT  124.36 275.98 250.08 276.66 ;
     RECT  261.66 275.64 282.74 277.85 ;
     RECT  261.66 277.85 282.28 278.36 ;
     RECT  6.6 276.35 18.94 278.7 ;
     RECT  261.66 278.36 278.14 278.7 ;
     RECT  261.66 278.7 277.68 279.21 ;
     RECT  30.97 232.8 32.51 280.345 ;
     RECT  58.11 191.66 59.65 280.345 ;
     RECT  71.68 275.98 113.93 280.345 ;
     RECT  248.09 276.66 250.08 280.345 ;
     RECT  42.48 268.7 46.08 281.42 ;
     RECT  71.68 280.345 104.26 281.42 ;
     RECT  71.68 281.42 103.8 281.76 ;
     RECT  124.36 276.66 236.06 281.76 ;
     RECT  261.66 279.21 277.22 281.93 ;
     RECT  71.68 281.76 103.34 281.96 ;
     RECT  10.28 278.7 18.94 283.065 ;
     RECT  44.54 281.42 46.08 283.065 ;
     RECT  125.96 281.76 236.06 283.065 ;
     RECT  261.66 281.93 274.46 283.065 ;
     RECT  10.28 283.065 11.34 288.66 ;
     RECT  64.56 281.96 103.34 288.66 ;
     RECT  129.88 283.065 227.54 288.66 ;
     RECT  248.56 280.345 250.08 288.66 ;
     RECT  271.56 283.065 274.46 288.66 ;
     RECT  132.18 288.66 133.7 288.73 ;
     RECT  249.02 288.66 250.08 288.73 ;
    LAYER met3 ;
     RECT  0.46 5.63 17.38 16.81 ;
     RECT  0.46 96.75 17.38 97.05 ;
     RECT  0.46 115.79 17.38 230.33 ;
     RECT  0.46 259.95 17.38 276.57 ;
     RECT  17.38 5.275 18.96 283.045 ;
     RECT  18.96 6.99 20.62 280.325 ;
     RECT  20.62 7.995 44.52 280.325 ;
     RECT  44.52 5.275 46.1 283.045 ;
     RECT  46.1 7.995 71.66 280.325 ;
     RECT  71.66 5.275 73.24 283.045 ;
     RECT  73.24 7.995 98.8 280.325 ;
     RECT  98.8 5.275 100.38 283.045 ;
     RECT  100.38 7.995 125.94 280.325 ;
     RECT  125.94 5.275 127.52 283.045 ;
     RECT  127.52 7.995 153.08 280.325 ;
     RECT  153.08 5.275 154.66 283.045 ;
     RECT  154.66 7.995 180.22 280.325 ;
     RECT  180.22 5.275 181.8 283.045 ;
     RECT  181.8 7.995 207.36 280.325 ;
     RECT  207.36 5.275 208.94 283.045 ;
     RECT  208.94 7.995 234.5 280.325 ;
     RECT  234.5 5.275 236.08 283.045 ;
     RECT  236.08 7.995 261.64 280.325 ;
     RECT  261.64 5.275 263.22 283.045 ;
     RECT  263.22 7.995 276.79 281.33 ;
     RECT  276.79 272.19 277 281.33 ;
     RECT  276.79 12.43 282.13 20.21 ;
     RECT  282.13 12.43 288.42 19.53 ;
     RECT  276.79 36.91 288.42 37.21 ;
     RECT  276.79 51.87 288.42 124.25 ;
     RECT  276.79 142.99 288.42 194.97 ;
     RECT  277 272.19 288.42 282.01 ;
     RECT  288.42 117.83 288.8 118.13 ;
    LAYER met4 ;
     RECT  17.37 5.2 18.97 7.92 ;
     RECT  44.51 5.2 46.11 7.92 ;
     RECT  71.65 5.2 73.25 7.92 ;
     RECT  98.79 5.2 100.39 7.92 ;
     RECT  125.93 5.2 127.53 7.92 ;
     RECT  153.07 5.2 154.67 7.92 ;
     RECT  180.21 5.2 181.81 7.92 ;
     RECT  207.35 5.2 208.95 7.92 ;
     RECT  234.49 5.2 236.09 7.92 ;
     RECT  261.63 5.2 263.23 7.92 ;
     RECT  17.37 7.92 276.8 280.4 ;
     RECT  17.37 280.4 18.97 283.12 ;
     RECT  44.51 280.4 46.11 283.12 ;
     RECT  71.65 280.4 73.25 283.12 ;
     RECT  98.79 280.4 100.39 283.12 ;
     RECT  125.93 280.4 127.53 283.12 ;
     RECT  153.07 280.4 154.67 283.12 ;
     RECT  180.21 280.4 181.81 283.12 ;
     RECT  207.35 280.4 208.95 283.12 ;
     RECT  234.49 280.4 236.09 283.12 ;
     RECT  261.63 280.4 263.23 283.12 ;
    LAYER met5 ;
     RECT  17.37 18.24 30.94 264.64 ;
     RECT  30.94 18.24 263.23 278.24 ;
     RECT  263.23 31.84 276.8 278.24 ;
  END
END serv_top
END LIBRARY
